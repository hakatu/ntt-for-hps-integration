library verilog;
use verilog.vl_types.all;
entity tb_barrett_reduction is
end tb_barrett_reduction;
