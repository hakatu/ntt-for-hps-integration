`timescale 1ns / 1ps 

////////////////////////////////////////////////////////////////////////////////// 

// Company:  

// Engineer:  

//  

// Create Date: 09/15/2023 04:17:28 PM 

// Design Name:  

// Module Name: wrap_tb 

// Project Name:  

// Target Devices:  

// Tool Versions:  

// Description:  

//  

// Dependencies:  

//  

// Revision: 

// Revision 0.01 - File Created 

// Additional Comments: 

//  

////////////////////////////////////////////////////////////////////////////////// 
`define SIMULATION
  

module wrap_tb_full; 

  
    reg aclr = 0;
	 
	 reg rd_req = 0;
	 
    reg clk = 0; 
    
    reg rst = 0; 
    
    reg start = 1;
    
    reg mode = 0; 
    
    reg we = 0;
    
    reg [7:0] address_ina;
    
    reg [7:0] address_inb;
    
    reg [15:0] data_ina;
    
    reg [15:0] data_inb;
    
    wire [15:0] data_out1;
    
    wire [15:0] data_out2;
    
    wire init_done;
    
    wire in_done;
    
    wire cal_done;
    
    wire done;
    
    wire wr_req;
	 
	 wire [31:0] rd_dat;
	 
	 wire rd_empty;
	 
	 wire [8:0] rd_used;
	 
	 wire wr_full;
	 
	 wire [8:0] wr_used;
	 
	 wire [31:0] temp;

//register to count the test number

reg [31:0] test_num;

  // Instantiate the wrap module 
	
//	wrap dut (
//		.clk(clk),
//		.rst(rst),
//		.start(start),
//		.mode(mode),
//		.we(we),
//		.address_ina(address_ina),
//		.address_inb(address_inb),
//		.data_ina(data_ina),
//		.data_inb(data_inb),
//		.data_out1(data_out1),
//		.data_out2(data_out2),
//		.init_done(init_done),
//		.in_done(in_done),
//		.cal_done(cal_done),
//		.done(done),
//		.wr_req(wr_req)
//		);

	wrap dut (
		.aclr(aclr),
		.rd_req(rd_req),
		.clk(clk),
		.rd_clk(clk),
		.rst(rst),
		.start(start),
		.mode(mode),
		.we(we),
		.address_ina(address_ina),
		.address_inb(address_inb),
		.data_ina(data_ina),
		.data_inb(data_inb),
		.data_out1(data_out1),
		.data_out2(data_out2),
		.init_done(init_done),
		.in_done(in_done),
		.cal_done(cal_done),
		.done(done),
		.wr_req(wr_req),
		.rd_dat(rd_dat),
		.rd_empty(rd_empty),
		.rd_used(rd_used),
		.wr_full(wr_full),
		.wr_used(wr_used),
		.temp(temp)
		);



  // Clock generation 

    always #5 clk = ~clk; 

  

  // Reset generation 

    initial begin 
test_num = 0;
			rst = 0;
			aclr = 1;
			#1000 
			aclr = 0;

/////Test Begin
////Begin test number #0//////////////
rst = 1;

//#1000
start = 1;
mode = 0; //NTT 0 // INTT 1

// Reset for a few clock cycles

#1000

rst = 0;
test_num = test_num + 1;
#1000
we = 1;
address_ina = 0;
address_inb = 1;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 2;
address_inb = 3;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 4;
address_inb = 5;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 6;
address_inb = 7;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 8;
address_inb = 9;
data_ina = 16'hffff;
data_inb = 16'hfffd;
#10;
address_ina = 10;
address_inb = 11;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 12;
address_inb = 13;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 14;
address_inb = 15;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 16;
address_inb = 17;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 18;
address_inb = 19;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 20;
address_inb = 21;
data_ina = 16'hfffe;
data_inb = 16'hffff;
#10;
address_ina = 22;
address_inb = 23;
data_ina = 16'hffff;
data_inb = 16'hfffe;
#10;
address_ina = 24;
address_inb = 25;
data_ina = 16'hfffd;
data_inb = 16'hffff;
#10;
address_ina = 26;
address_inb = 27;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 28;
address_inb = 29;
data_ina = 16'h0;
data_inb = 16'h3;
#10;
address_ina = 30;
address_inb = 31;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 32;
address_inb = 33;
data_ina = 16'hfffe;
data_inb = 16'h1;
#10;
address_ina = 34;
address_inb = 35;
data_ina = 16'hfffe;
data_inb = 16'hffff;
#10;
address_ina = 36;
address_inb = 37;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 38;
address_inb = 39;
data_ina = 16'h2;
data_inb = 16'hffff;
#10;
address_ina = 40;
address_inb = 41;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 42;
address_inb = 43;
data_ina = 16'hffff;
data_inb = 16'hfffe;
#10;
address_ina = 44;
address_inb = 45;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 46;
address_inb = 47;
data_ina = 16'h2;
data_inb = 16'h2;
#10;
address_ina = 48;
address_inb = 49;
data_ina = 16'hffff;
data_inb = 16'h3;
#10;
address_ina = 50;
address_inb = 51;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 52;
address_inb = 53;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 54;
address_inb = 55;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 56;
address_inb = 57;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 58;
address_inb = 59;
data_ina = 16'h0;
data_inb = 16'h2;
#10;
address_ina = 60;
address_inb = 61;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 62;
address_inb = 63;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 64;
address_inb = 65;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 66;
address_inb = 67;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 68;
address_inb = 69;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 70;
address_inb = 71;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 72;
address_inb = 73;
data_ina = 16'hffff;
data_inb = 16'h2;
#10;
address_ina = 74;
address_inb = 75;
data_ina = 16'h0;
data_inb = 16'hfffe;
#10;
address_ina = 76;
address_inb = 77;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 78;
address_inb = 79;
data_ina = 16'h2;
data_inb = 16'h0;
#10;
address_ina = 80;
address_inb = 81;
data_ina = 16'h2;
data_inb = 16'h1;
#10;
address_ina = 82;
address_inb = 83;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 84;
address_inb = 85;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 86;
address_inb = 87;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 88;
address_inb = 89;
data_ina = 16'h1;
data_inb = 16'hfffd;
#10;
address_ina = 90;
address_inb = 91;
data_ina = 16'h2;
data_inb = 16'h0;
#10;
address_ina = 92;
address_inb = 93;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 94;
address_inb = 95;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 96;
address_inb = 97;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 98;
address_inb = 99;
data_ina = 16'h0;
data_inb = 16'h2;
#10;
address_ina = 100;
address_inb = 101;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 102;
address_inb = 103;
data_ina = 16'hfffe;
data_inb = 16'h0;
#10;
address_ina = 104;
address_inb = 105;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 106;
address_inb = 107;
data_ina = 16'h3;
data_inb = 16'h0;
#10;
address_ina = 108;
address_inb = 109;
data_ina = 16'h2;
data_inb = 16'h1;
#10;
address_ina = 110;
address_inb = 111;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 112;
address_inb = 113;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 114;
address_inb = 115;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 116;
address_inb = 117;
data_ina = 16'h1;
data_inb = 16'hfffe;
#10;
address_ina = 118;
address_inb = 119;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 120;
address_inb = 121;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 122;
address_inb = 123;
data_ina = 16'hffff;
data_inb = 16'hfffe;
#10;
address_ina = 124;
address_inb = 125;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 126;
address_inb = 127;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 128;
address_inb = 129;
data_ina = 16'h0;
data_inb = 16'h3;
#10;
address_ina = 130;
address_inb = 131;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 132;
address_inb = 133;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 134;
address_inb = 135;
data_ina = 16'hfffe;
data_inb = 16'h0;
#10;
address_ina = 136;
address_inb = 137;
data_ina = 16'h1;
data_inb = 16'hfffe;
#10;
address_ina = 138;
address_inb = 139;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 140;
address_inb = 141;
data_ina = 16'h1;
data_inb = 16'h2;
#10;
address_ina = 142;
address_inb = 143;
data_ina = 16'h2;
data_inb = 16'h0;
#10;
address_ina = 144;
address_inb = 145;
data_ina = 16'hfffe;
data_inb = 16'h0;
#10;
address_ina = 146;
address_inb = 147;
data_ina = 16'h0;
data_inb = 16'hfffd;
#10;
address_ina = 148;
address_inb = 149;
data_ina = 16'hfffd;
data_inb = 16'h1;
#10;
address_ina = 150;
address_inb = 151;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 152;
address_inb = 153;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 154;
address_inb = 155;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 156;
address_inb = 157;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 158;
address_inb = 159;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 160;
address_inb = 161;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 162;
address_inb = 163;
data_ina = 16'hfffd;
data_inb = 16'h0;
#10;
address_ina = 164;
address_inb = 165;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 166;
address_inb = 167;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 168;
address_inb = 169;
data_ina = 16'hfffe;
data_inb = 16'h0;
#10;
address_ina = 170;
address_inb = 171;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 172;
address_inb = 173;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 174;
address_inb = 175;
data_ina = 16'hffff;
data_inb = 16'h2;
#10;
address_ina = 176;
address_inb = 177;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 178;
address_inb = 179;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 180;
address_inb = 181;
data_ina = 16'hfffe;
data_inb = 16'h0;
#10;
address_ina = 182;
address_inb = 183;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 184;
address_inb = 185;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 186;
address_inb = 187;
data_ina = 16'hffff;
data_inb = 16'h2;
#10;
address_ina = 188;
address_inb = 189;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 190;
address_inb = 191;
data_ina = 16'h2;
data_inb = 16'h0;
#10;
address_ina = 192;
address_inb = 193;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 194;
address_inb = 195;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 196;
address_inb = 197;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 198;
address_inb = 199;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 200;
address_inb = 201;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 202;
address_inb = 203;
data_ina = 16'h2;
data_inb = 16'h1;
#10;
address_ina = 204;
address_inb = 205;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 206;
address_inb = 207;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 208;
address_inb = 209;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 210;
address_inb = 211;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 212;
address_inb = 213;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 214;
address_inb = 215;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 216;
address_inb = 217;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 218;
address_inb = 219;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 220;
address_inb = 221;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 222;
address_inb = 223;
data_ina = 16'hfffe;
data_inb = 16'h1;
#10;
address_ina = 224;
address_inb = 225;
data_ina = 16'hfffe;
data_inb = 16'h1;
#10;
address_ina = 226;
address_inb = 227;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 228;
address_inb = 229;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 230;
address_inb = 231;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 232;
address_inb = 233;
data_ina = 16'hfffe;
data_inb = 16'h1;
#10;
address_ina = 234;
address_inb = 235;
data_ina = 16'hfffd;
data_inb = 16'h1;
#10;
address_ina = 236;
address_inb = 237;
data_ina = 16'h2;
data_inb = 16'h2;
#10;
address_ina = 238;
address_inb = 239;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 240;
address_inb = 241;
data_ina = 16'hfffe;
data_inb = 16'hffff;
#10;
address_ina = 242;
address_inb = 243;
data_ina = 16'h0;
data_inb = 16'hfffe;
#10;
address_ina = 244;
address_inb = 245;
data_ina = 16'h2;
data_inb = 16'h0;
#10;
address_ina = 246;
address_inb = 247;
data_ina = 16'hfffe;
data_inb = 16'h2;
#10;
address_ina = 248;
address_inb = 249;
data_ina = 16'h1;
data_inb = 16'h2;
#10;
address_ina = 250;
address_inb = 251;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 252;
address_inb = 253;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 254;
address_inb = 255;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
        wait(init_done);
        #30
        we = 0;
        // Start processing
         
		  #38000

        start = 0;



//        wait (wr_req);
//		  wait (!wr_req);
//		   rd_req = 1;
		  wait(done);
		  #20000
rd_req = 1;
        #70 
		  start = 1;
		 #80 
wait(rd_empty)
rd_req = 0;

$display("Finished the NTT test Number %d",test_num);
////Begin test number #1//////////////
rst = 1;

//#1000
start = 1;
mode = 0; //NTT 0 // INTT 1

// Reset for a few clock cycles

#1000

rst = 0;
test_num = test_num + 1;
#1000
we = 1;
address_ina = 0;
address_inb = 1;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 2;
address_inb = 3;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 4;
address_inb = 5;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 6;
address_inb = 7;
data_ina = 16'hfffe;
data_inb = 16'h1;
#10;
address_ina = 8;
address_inb = 9;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 10;
address_inb = 11;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 12;
address_inb = 13;
data_ina = 16'hfffe;
data_inb = 16'hffff;
#10;
address_ina = 14;
address_inb = 15;
data_ina = 16'hfffe;
data_inb = 16'hffff;
#10;
address_ina = 16;
address_inb = 17;
data_ina = 16'h3;
data_inb = 16'h0;
#10;
address_ina = 18;
address_inb = 19;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 20;
address_inb = 21;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 22;
address_inb = 23;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 24;
address_inb = 25;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 26;
address_inb = 27;
data_ina = 16'hffff;
data_inb = 16'hfffe;
#10;
address_ina = 28;
address_inb = 29;
data_ina = 16'h2;
data_inb = 16'hfffe;
#10;
address_ina = 30;
address_inb = 31;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 32;
address_inb = 33;
data_ina = 16'h2;
data_inb = 16'h2;
#10;
address_ina = 34;
address_inb = 35;
data_ina = 16'hfffe;
data_inb = 16'h0;
#10;
address_ina = 36;
address_inb = 37;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 38;
address_inb = 39;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 40;
address_inb = 41;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 42;
address_inb = 43;
data_ina = 16'h2;
data_inb = 16'hffff;
#10;
address_ina = 44;
address_inb = 45;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 46;
address_inb = 47;
data_ina = 16'hffff;
data_inb = 16'hfffe;
#10;
address_ina = 48;
address_inb = 49;
data_ina = 16'hfffe;
data_inb = 16'h0;
#10;
address_ina = 50;
address_inb = 51;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 52;
address_inb = 53;
data_ina = 16'h3;
data_inb = 16'h0;
#10;
address_ina = 54;
address_inb = 55;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 56;
address_inb = 57;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 58;
address_inb = 59;
data_ina = 16'h2;
data_inb = 16'h1;
#10;
address_ina = 60;
address_inb = 61;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 62;
address_inb = 63;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 64;
address_inb = 65;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 66;
address_inb = 67;
data_ina = 16'hfffe;
data_inb = 16'h0;
#10;
address_ina = 68;
address_inb = 69;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 70;
address_inb = 71;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 72;
address_inb = 73;
data_ina = 16'h0;
data_inb = 16'h2;
#10;
address_ina = 74;
address_inb = 75;
data_ina = 16'hffff;
data_inb = 16'h2;
#10;
address_ina = 76;
address_inb = 77;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 78;
address_inb = 79;
data_ina = 16'hffff;
data_inb = 16'hfffe;
#10;
address_ina = 80;
address_inb = 81;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 82;
address_inb = 83;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 84;
address_inb = 85;
data_ina = 16'hffff;
data_inb = 16'h3;
#10;
address_ina = 86;
address_inb = 87;
data_ina = 16'h2;
data_inb = 16'hfffe;
#10;
address_ina = 88;
address_inb = 89;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 90;
address_inb = 91;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 92;
address_inb = 93;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 94;
address_inb = 95;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 96;
address_inb = 97;
data_ina = 16'h0;
data_inb = 16'hfffe;
#10;
address_ina = 98;
address_inb = 99;
data_ina = 16'hfffe;
data_inb = 16'h1;
#10;
address_ina = 100;
address_inb = 101;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 102;
address_inb = 103;
data_ina = 16'hfffe;
data_inb = 16'hffff;
#10;
address_ina = 104;
address_inb = 105;
data_ina = 16'hfffe;
data_inb = 16'hffff;
#10;
address_ina = 106;
address_inb = 107;
data_ina = 16'h2;
data_inb = 16'hffff;
#10;
address_ina = 108;
address_inb = 109;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 110;
address_inb = 111;
data_ina = 16'h0;
data_inb = 16'h2;
#10;
address_ina = 112;
address_inb = 113;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 114;
address_inb = 115;
data_ina = 16'h2;
data_inb = 16'h0;
#10;
address_ina = 116;
address_inb = 117;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 118;
address_inb = 119;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 120;
address_inb = 121;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 122;
address_inb = 123;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 124;
address_inb = 125;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 126;
address_inb = 127;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 128;
address_inb = 129;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 130;
address_inb = 131;
data_ina = 16'h2;
data_inb = 16'h1;
#10;
address_ina = 132;
address_inb = 133;
data_ina = 16'h2;
data_inb = 16'h1;
#10;
address_ina = 134;
address_inb = 135;
data_ina = 16'h2;
data_inb = 16'h1;
#10;
address_ina = 136;
address_inb = 137;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 138;
address_inb = 139;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 140;
address_inb = 141;
data_ina = 16'h2;
data_inb = 16'hffff;
#10;
address_ina = 142;
address_inb = 143;
data_ina = 16'hfffe;
data_inb = 16'h0;
#10;
address_ina = 144;
address_inb = 145;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 146;
address_inb = 147;
data_ina = 16'h1;
data_inb = 16'h2;
#10;
address_ina = 148;
address_inb = 149;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 150;
address_inb = 151;
data_ina = 16'h2;
data_inb = 16'hffff;
#10;
address_ina = 152;
address_inb = 153;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 154;
address_inb = 155;
data_ina = 16'hffff;
data_inb = 16'h2;
#10;
address_ina = 156;
address_inb = 157;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 158;
address_inb = 159;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 160;
address_inb = 161;
data_ina = 16'hffff;
data_inb = 16'h2;
#10;
address_ina = 162;
address_inb = 163;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 164;
address_inb = 165;
data_ina = 16'h0;
data_inb = 16'hfffe;
#10;
address_ina = 166;
address_inb = 167;
data_ina = 16'h1;
data_inb = 16'h2;
#10;
address_ina = 168;
address_inb = 169;
data_ina = 16'h2;
data_inb = 16'h0;
#10;
address_ina = 170;
address_inb = 171;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 172;
address_inb = 173;
data_ina = 16'hffff;
data_inb = 16'h2;
#10;
address_ina = 174;
address_inb = 175;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 176;
address_inb = 177;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 178;
address_inb = 179;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 180;
address_inb = 181;
data_ina = 16'h2;
data_inb = 16'h0;
#10;
address_ina = 182;
address_inb = 183;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 184;
address_inb = 185;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 186;
address_inb = 187;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 188;
address_inb = 189;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 190;
address_inb = 191;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 192;
address_inb = 193;
data_ina = 16'h0;
data_inb = 16'hfffe;
#10;
address_ina = 194;
address_inb = 195;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 196;
address_inb = 197;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 198;
address_inb = 199;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 200;
address_inb = 201;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 202;
address_inb = 203;
data_ina = 16'hffff;
data_inb = 16'h2;
#10;
address_ina = 204;
address_inb = 205;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 206;
address_inb = 207;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 208;
address_inb = 209;
data_ina = 16'hfffe;
data_inb = 16'h1;
#10;
address_ina = 210;
address_inb = 211;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 212;
address_inb = 213;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 214;
address_inb = 215;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 216;
address_inb = 217;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 218;
address_inb = 219;
data_ina = 16'hfffe;
data_inb = 16'hffff;
#10;
address_ina = 220;
address_inb = 221;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 222;
address_inb = 223;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 224;
address_inb = 225;
data_ina = 16'h0;
data_inb = 16'h2;
#10;
address_ina = 226;
address_inb = 227;
data_ina = 16'h2;
data_inb = 16'hfffd;
#10;
address_ina = 228;
address_inb = 229;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 230;
address_inb = 231;
data_ina = 16'h2;
data_inb = 16'h1;
#10;
address_ina = 232;
address_inb = 233;
data_ina = 16'hfffe;
data_inb = 16'h0;
#10;
address_ina = 234;
address_inb = 235;
data_ina = 16'hfffe;
data_inb = 16'hfffe;
#10;
address_ina = 236;
address_inb = 237;
data_ina = 16'h2;
data_inb = 16'h0;
#10;
address_ina = 238;
address_inb = 239;
data_ina = 16'hfffe;
data_inb = 16'h1;
#10;
address_ina = 240;
address_inb = 241;
data_ina = 16'hffff;
data_inb = 16'h2;
#10;
address_ina = 242;
address_inb = 243;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 244;
address_inb = 245;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 246;
address_inb = 247;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 248;
address_inb = 249;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 250;
address_inb = 251;
data_ina = 16'h0;
data_inb = 16'hfffe;
#10;
address_ina = 252;
address_inb = 253;
data_ina = 16'h3;
data_inb = 16'h2;
#10;
address_ina = 254;
address_inb = 255;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
        wait(init_done);
        #30
        we = 0;
        // Start processing
         
		  #38000

        start = 0;



//        wait (wr_req);
//		  wait (!wr_req);
//		   rd_req = 1;
		  wait(done);
		  #20000
rd_req = 1;
        #70 
		  start = 1;
		 #80 
wait(rd_empty)
rd_req = 0;

$display("Finished the NTT test Number %d",test_num);
////Begin test number #2//////////////
rst = 1;

//#1000
start = 1;
mode = 0; //NTT 0 // INTT 1

// Reset for a few clock cycles

#1000

rst = 0;
test_num = test_num + 1;
#1000
we = 1;
address_ina = 0;
address_inb = 1;
data_ina = 16'hfffe;
data_inb = 16'h1;
#10;
address_ina = 2;
address_inb = 3;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 4;
address_inb = 5;
data_ina = 16'h2;
data_inb = 16'h0;
#10;
address_ina = 6;
address_inb = 7;
data_ina = 16'h1;
data_inb = 16'h2;
#10;
address_ina = 8;
address_inb = 9;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 10;
address_inb = 11;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 12;
address_inb = 13;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 14;
address_inb = 15;
data_ina = 16'hfffd;
data_inb = 16'hffff;
#10;
address_ina = 16;
address_inb = 17;
data_ina = 16'h0;
data_inb = 16'h2;
#10;
address_ina = 18;
address_inb = 19;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 20;
address_inb = 21;
data_ina = 16'h0;
data_inb = 16'hfffd;
#10;
address_ina = 22;
address_inb = 23;
data_ina = 16'h2;
data_inb = 16'h1;
#10;
address_ina = 24;
address_inb = 25;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 26;
address_inb = 27;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 28;
address_inb = 29;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 30;
address_inb = 31;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 32;
address_inb = 33;
data_ina = 16'h3;
data_inb = 16'h0;
#10;
address_ina = 34;
address_inb = 35;
data_ina = 16'h2;
data_inb = 16'h0;
#10;
address_ina = 36;
address_inb = 37;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 38;
address_inb = 39;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 40;
address_inb = 41;
data_ina = 16'h1;
data_inb = 16'hfffd;
#10;
address_ina = 42;
address_inb = 43;
data_ina = 16'hfffe;
data_inb = 16'h1;
#10;
address_ina = 44;
address_inb = 45;
data_ina = 16'h2;
data_inb = 16'hffff;
#10;
address_ina = 46;
address_inb = 47;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 48;
address_inb = 49;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 50;
address_inb = 51;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 52;
address_inb = 53;
data_ina = 16'h1;
data_inb = 16'hfffe;
#10;
address_ina = 54;
address_inb = 55;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 56;
address_inb = 57;
data_ina = 16'hfffd;
data_inb = 16'h0;
#10;
address_ina = 58;
address_inb = 59;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 60;
address_inb = 61;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 62;
address_inb = 63;
data_ina = 16'hffff;
data_inb = 16'hfffe;
#10;
address_ina = 64;
address_inb = 65;
data_ina = 16'h3;
data_inb = 16'h1;
#10;
address_ina = 66;
address_inb = 67;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 68;
address_inb = 69;
data_ina = 16'h0;
data_inb = 16'h3;
#10;
address_ina = 70;
address_inb = 71;
data_ina = 16'h0;
data_inb = 16'hfffd;
#10;
address_ina = 72;
address_inb = 73;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 74;
address_inb = 75;
data_ina = 16'h2;
data_inb = 16'h1;
#10;
address_ina = 76;
address_inb = 77;
data_ina = 16'h2;
data_inb = 16'h2;
#10;
address_ina = 78;
address_inb = 79;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 80;
address_inb = 81;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 82;
address_inb = 83;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 84;
address_inb = 85;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 86;
address_inb = 87;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 88;
address_inb = 89;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 90;
address_inb = 91;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 92;
address_inb = 93;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 94;
address_inb = 95;
data_ina = 16'hfffe;
data_inb = 16'h1;
#10;
address_ina = 96;
address_inb = 97;
data_ina = 16'hfffe;
data_inb = 16'h0;
#10;
address_ina = 98;
address_inb = 99;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 100;
address_inb = 101;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 102;
address_inb = 103;
data_ina = 16'h2;
data_inb = 16'h0;
#10;
address_ina = 104;
address_inb = 105;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 106;
address_inb = 107;
data_ina = 16'h1;
data_inb = 16'hfffe;
#10;
address_ina = 108;
address_inb = 109;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 110;
address_inb = 111;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 112;
address_inb = 113;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 114;
address_inb = 115;
data_ina = 16'hfffe;
data_inb = 16'hfffe;
#10;
address_ina = 116;
address_inb = 117;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 118;
address_inb = 119;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 120;
address_inb = 121;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 122;
address_inb = 123;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 124;
address_inb = 125;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 126;
address_inb = 127;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 128;
address_inb = 129;
data_ina = 16'h1;
data_inb = 16'hfffe;
#10;
address_ina = 130;
address_inb = 131;
data_ina = 16'h1;
data_inb = 16'h2;
#10;
address_ina = 132;
address_inb = 133;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 134;
address_inb = 135;
data_ina = 16'h2;
data_inb = 16'h1;
#10;
address_ina = 136;
address_inb = 137;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 138;
address_inb = 139;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 140;
address_inb = 141;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 142;
address_inb = 143;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 144;
address_inb = 145;
data_ina = 16'h2;
data_inb = 16'h2;
#10;
address_ina = 146;
address_inb = 147;
data_ina = 16'h0;
data_inb = 16'hfffe;
#10;
address_ina = 148;
address_inb = 149;
data_ina = 16'hffff;
data_inb = 16'h2;
#10;
address_ina = 150;
address_inb = 151;
data_ina = 16'h0;
data_inb = 16'hfffe;
#10;
address_ina = 152;
address_inb = 153;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 154;
address_inb = 155;
data_ina = 16'h0;
data_inb = 16'hfffe;
#10;
address_ina = 156;
address_inb = 157;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 158;
address_inb = 159;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 160;
address_inb = 161;
data_ina = 16'h0;
data_inb = 16'hfffe;
#10;
address_ina = 162;
address_inb = 163;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 164;
address_inb = 165;
data_ina = 16'h2;
data_inb = 16'hffff;
#10;
address_ina = 166;
address_inb = 167;
data_ina = 16'hfffe;
data_inb = 16'h1;
#10;
address_ina = 168;
address_inb = 169;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 170;
address_inb = 171;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 172;
address_inb = 173;
data_ina = 16'h0;
data_inb = 16'h2;
#10;
address_ina = 174;
address_inb = 175;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 176;
address_inb = 177;
data_ina = 16'h2;
data_inb = 16'hffff;
#10;
address_ina = 178;
address_inb = 179;
data_ina = 16'hffff;
data_inb = 16'h2;
#10;
address_ina = 180;
address_inb = 181;
data_ina = 16'h0;
data_inb = 16'h2;
#10;
address_ina = 182;
address_inb = 183;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 184;
address_inb = 185;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 186;
address_inb = 187;
data_ina = 16'hffff;
data_inb = 16'h2;
#10;
address_ina = 188;
address_inb = 189;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 190;
address_inb = 191;
data_ina = 16'h2;
data_inb = 16'h1;
#10;
address_ina = 192;
address_inb = 193;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 194;
address_inb = 195;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 196;
address_inb = 197;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 198;
address_inb = 199;
data_ina = 16'h0;
data_inb = 16'hfffe;
#10;
address_ina = 200;
address_inb = 201;
data_ina = 16'h2;
data_inb = 16'hfffd;
#10;
address_ina = 202;
address_inb = 203;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 204;
address_inb = 205;
data_ina = 16'h1;
data_inb = 16'h2;
#10;
address_ina = 206;
address_inb = 207;
data_ina = 16'h1;
data_inb = 16'h2;
#10;
address_ina = 208;
address_inb = 209;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 210;
address_inb = 211;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 212;
address_inb = 213;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 214;
address_inb = 215;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 216;
address_inb = 217;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 218;
address_inb = 219;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 220;
address_inb = 221;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 222;
address_inb = 223;
data_ina = 16'h0;
data_inb = 16'hfffe;
#10;
address_ina = 224;
address_inb = 225;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 226;
address_inb = 227;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 228;
address_inb = 229;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 230;
address_inb = 231;
data_ina = 16'h0;
data_inb = 16'hfffe;
#10;
address_ina = 232;
address_inb = 233;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 234;
address_inb = 235;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 236;
address_inb = 237;
data_ina = 16'hffff;
data_inb = 16'h2;
#10;
address_ina = 238;
address_inb = 239;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 240;
address_inb = 241;
data_ina = 16'h3;
data_inb = 16'h1;
#10;
address_ina = 242;
address_inb = 243;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 244;
address_inb = 245;
data_ina = 16'h2;
data_inb = 16'hffff;
#10;
address_ina = 246;
address_inb = 247;
data_ina = 16'hfffe;
data_inb = 16'hffff;
#10;
address_ina = 248;
address_inb = 249;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 250;
address_inb = 251;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 252;
address_inb = 253;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 254;
address_inb = 255;
data_ina = 16'hfffe;
data_inb = 16'h0;
#10;
        wait(init_done);
        #30
        we = 0;
        // Start processing
         
		  #38000

        start = 0;



//        wait (wr_req);
//		  wait (!wr_req);
//		   rd_req = 1;
		  wait(done);
		  #20000
rd_req = 1;
        #70 
		  start = 1;
		 #80 
wait(rd_empty)
rd_req = 0;

$display("Finished the NTT test Number %d",test_num);
////Begin test number #3//////////////
rst = 1;

//#1000
start = 1;
mode = 0; //NTT 0 // INTT 1

// Reset for a few clock cycles

#1000

rst = 0;
test_num = test_num + 1;
#1000
we = 1;
address_ina = 0;
address_inb = 1;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 2;
address_inb = 3;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 4;
address_inb = 5;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 6;
address_inb = 7;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 8;
address_inb = 9;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 10;
address_inb = 11;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 12;
address_inb = 13;
data_ina = 16'h2;
data_inb = 16'h0;
#10;
address_ina = 14;
address_inb = 15;
data_ina = 16'h2;
data_inb = 16'h0;
#10;
address_ina = 16;
address_inb = 17;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 18;
address_inb = 19;
data_ina = 16'hfffe;
data_inb = 16'hffff;
#10;
address_ina = 20;
address_inb = 21;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 22;
address_inb = 23;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 24;
address_inb = 25;
data_ina = 16'hfffe;
data_inb = 16'hffff;
#10;
address_ina = 26;
address_inb = 27;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 28;
address_inb = 29;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 30;
address_inb = 31;
data_ina = 16'h2;
data_inb = 16'hfffe;
#10;
address_ina = 32;
address_inb = 33;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 34;
address_inb = 35;
data_ina = 16'hfffd;
data_inb = 16'h1;
#10;
address_ina = 36;
address_inb = 37;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 38;
address_inb = 39;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 40;
address_inb = 41;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 42;
address_inb = 43;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 44;
address_inb = 45;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 46;
address_inb = 47;
data_ina = 16'h2;
data_inb = 16'h0;
#10;
address_ina = 48;
address_inb = 49;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 50;
address_inb = 51;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 52;
address_inb = 53;
data_ina = 16'h2;
data_inb = 16'hfffe;
#10;
address_ina = 54;
address_inb = 55;
data_ina = 16'hfffe;
data_inb = 16'h1;
#10;
address_ina = 56;
address_inb = 57;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 58;
address_inb = 59;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 60;
address_inb = 61;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 62;
address_inb = 63;
data_ina = 16'hfffe;
data_inb = 16'hfffe;
#10;
address_ina = 64;
address_inb = 65;
data_ina = 16'h2;
data_inb = 16'h2;
#10;
address_ina = 66;
address_inb = 67;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 68;
address_inb = 69;
data_ina = 16'hfffe;
data_inb = 16'hffff;
#10;
address_ina = 70;
address_inb = 71;
data_ina = 16'h0;
data_inb = 16'hfffe;
#10;
address_ina = 72;
address_inb = 73;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 74;
address_inb = 75;
data_ina = 16'h1;
data_inb = 16'h2;
#10;
address_ina = 76;
address_inb = 77;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 78;
address_inb = 79;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 80;
address_inb = 81;
data_ina = 16'hffff;
data_inb = 16'hfffe;
#10;
address_ina = 82;
address_inb = 83;
data_ina = 16'h0;
data_inb = 16'h2;
#10;
address_ina = 84;
address_inb = 85;
data_ina = 16'h1;
data_inb = 16'hfffe;
#10;
address_ina = 86;
address_inb = 87;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 88;
address_inb = 89;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 90;
address_inb = 91;
data_ina = 16'hfffe;
data_inb = 16'h0;
#10;
address_ina = 92;
address_inb = 93;
data_ina = 16'h2;
data_inb = 16'h2;
#10;
address_ina = 94;
address_inb = 95;
data_ina = 16'h1;
data_inb = 16'hfffe;
#10;
address_ina = 96;
address_inb = 97;
data_ina = 16'h0;
data_inb = 16'hfffd;
#10;
address_ina = 98;
address_inb = 99;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 100;
address_inb = 101;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 102;
address_inb = 103;
data_ina = 16'h0;
data_inb = 16'h2;
#10;
address_ina = 104;
address_inb = 105;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 106;
address_inb = 107;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 108;
address_inb = 109;
data_ina = 16'h0;
data_inb = 16'h2;
#10;
address_ina = 110;
address_inb = 111;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 112;
address_inb = 113;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 114;
address_inb = 115;
data_ina = 16'h0;
data_inb = 16'h2;
#10;
address_ina = 116;
address_inb = 117;
data_ina = 16'hfffe;
data_inb = 16'h0;
#10;
address_ina = 118;
address_inb = 119;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 120;
address_inb = 121;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 122;
address_inb = 123;
data_ina = 16'h0;
data_inb = 16'h2;
#10;
address_ina = 124;
address_inb = 125;
data_ina = 16'hfffe;
data_inb = 16'hfffe;
#10;
address_ina = 126;
address_inb = 127;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 128;
address_inb = 129;
data_ina = 16'hfffe;
data_inb = 16'h2;
#10;
address_ina = 130;
address_inb = 131;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 132;
address_inb = 133;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 134;
address_inb = 135;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 136;
address_inb = 137;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 138;
address_inb = 139;
data_ina = 16'h2;
data_inb = 16'h0;
#10;
address_ina = 140;
address_inb = 141;
data_ina = 16'h2;
data_inb = 16'h2;
#10;
address_ina = 142;
address_inb = 143;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 144;
address_inb = 145;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 146;
address_inb = 147;
data_ina = 16'hfffd;
data_inb = 16'h0;
#10;
address_ina = 148;
address_inb = 149;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 150;
address_inb = 151;
data_ina = 16'h0;
data_inb = 16'h2;
#10;
address_ina = 152;
address_inb = 153;
data_ina = 16'h2;
data_inb = 16'h0;
#10;
address_ina = 154;
address_inb = 155;
data_ina = 16'h3;
data_inb = 16'hfffd;
#10;
address_ina = 156;
address_inb = 157;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 158;
address_inb = 159;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 160;
address_inb = 161;
data_ina = 16'hfffe;
data_inb = 16'h0;
#10;
address_ina = 162;
address_inb = 163;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 164;
address_inb = 165;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 166;
address_inb = 167;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 168;
address_inb = 169;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 170;
address_inb = 171;
data_ina = 16'hffff;
data_inb = 16'hfffe;
#10;
address_ina = 172;
address_inb = 173;
data_ina = 16'h2;
data_inb = 16'hffff;
#10;
address_ina = 174;
address_inb = 175;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 176;
address_inb = 177;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 178;
address_inb = 179;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 180;
address_inb = 181;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 182;
address_inb = 183;
data_ina = 16'h0;
data_inb = 16'hfffe;
#10;
address_ina = 184;
address_inb = 185;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 186;
address_inb = 187;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 188;
address_inb = 189;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 190;
address_inb = 191;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 192;
address_inb = 193;
data_ina = 16'hfffe;
data_inb = 16'h0;
#10;
address_ina = 194;
address_inb = 195;
data_ina = 16'hffff;
data_inb = 16'h2;
#10;
address_ina = 196;
address_inb = 197;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 198;
address_inb = 199;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 200;
address_inb = 201;
data_ina = 16'hfffe;
data_inb = 16'h0;
#10;
address_ina = 202;
address_inb = 203;
data_ina = 16'hfffe;
data_inb = 16'h1;
#10;
address_ina = 204;
address_inb = 205;
data_ina = 16'h2;
data_inb = 16'h1;
#10;
address_ina = 206;
address_inb = 207;
data_ina = 16'h3;
data_inb = 16'h1;
#10;
address_ina = 208;
address_inb = 209;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 210;
address_inb = 211;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 212;
address_inb = 213;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 214;
address_inb = 215;
data_ina = 16'h1;
data_inb = 16'hfffe;
#10;
address_ina = 216;
address_inb = 217;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 218;
address_inb = 219;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 220;
address_inb = 221;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 222;
address_inb = 223;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 224;
address_inb = 225;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 226;
address_inb = 227;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 228;
address_inb = 229;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 230;
address_inb = 231;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 232;
address_inb = 233;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 234;
address_inb = 235;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 236;
address_inb = 237;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 238;
address_inb = 239;
data_ina = 16'h2;
data_inb = 16'hffff;
#10;
address_ina = 240;
address_inb = 241;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 242;
address_inb = 243;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 244;
address_inb = 245;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 246;
address_inb = 247;
data_ina = 16'h2;
data_inb = 16'hffff;
#10;
address_ina = 248;
address_inb = 249;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 250;
address_inb = 251;
data_ina = 16'h2;
data_inb = 16'h2;
#10;
address_ina = 252;
address_inb = 253;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 254;
address_inb = 255;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
        wait(init_done);
        #30
        we = 0;
        // Start processing
         
		  #38000

        start = 0;



//        wait (wr_req);
//		  wait (!wr_req);
//		   rd_req = 1;
		  wait(done);
		  #20000
rd_req = 1;
        #70 
		  start = 1;
		 #80 
wait(rd_empty)
rd_req = 0;

$display("Finished the NTT test Number %d",test_num);
////Begin test number #4//////////////
rst = 1;

//#1000
start = 1;
mode = 0; //NTT 0 // INTT 1

// Reset for a few clock cycles

#1000

rst = 0;
test_num = test_num + 1;
#1000
we = 1;
address_ina = 0;
address_inb = 1;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 2;
address_inb = 3;
data_ina = 16'h2;
data_inb = 16'hffff;
#10;
address_ina = 4;
address_inb = 5;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 6;
address_inb = 7;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 8;
address_inb = 9;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 10;
address_inb = 11;
data_ina = 16'hfffe;
data_inb = 16'h1;
#10;
address_ina = 12;
address_inb = 13;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 14;
address_inb = 15;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 16;
address_inb = 17;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 18;
address_inb = 19;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 20;
address_inb = 21;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 22;
address_inb = 23;
data_ina = 16'h0;
data_inb = 16'h2;
#10;
address_ina = 24;
address_inb = 25;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 26;
address_inb = 27;
data_ina = 16'h0;
data_inb = 16'h2;
#10;
address_ina = 28;
address_inb = 29;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 30;
address_inb = 31;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 32;
address_inb = 33;
data_ina = 16'hfffe;
data_inb = 16'hfffd;
#10;
address_ina = 34;
address_inb = 35;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 36;
address_inb = 37;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 38;
address_inb = 39;
data_ina = 16'h1;
data_inb = 16'h2;
#10;
address_ina = 40;
address_inb = 41;
data_ina = 16'h2;
data_inb = 16'h0;
#10;
address_ina = 42;
address_inb = 43;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 44;
address_inb = 45;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 46;
address_inb = 47;
data_ina = 16'h2;
data_inb = 16'hffff;
#10;
address_ina = 48;
address_inb = 49;
data_ina = 16'hfffd;
data_inb = 16'h2;
#10;
address_ina = 50;
address_inb = 51;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 52;
address_inb = 53;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 54;
address_inb = 55;
data_ina = 16'h0;
data_inb = 16'hfffe;
#10;
address_ina = 56;
address_inb = 57;
data_ina = 16'hfffe;
data_inb = 16'h0;
#10;
address_ina = 58;
address_inb = 59;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 60;
address_inb = 61;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 62;
address_inb = 63;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 64;
address_inb = 65;
data_ina = 16'hfffe;
data_inb = 16'h1;
#10;
address_ina = 66;
address_inb = 67;
data_ina = 16'hfffe;
data_inb = 16'h0;
#10;
address_ina = 68;
address_inb = 69;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 70;
address_inb = 71;
data_ina = 16'h2;
data_inb = 16'h1;
#10;
address_ina = 72;
address_inb = 73;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 74;
address_inb = 75;
data_ina = 16'h2;
data_inb = 16'h0;
#10;
address_ina = 76;
address_inb = 77;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 78;
address_inb = 79;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 80;
address_inb = 81;
data_ina = 16'hffff;
data_inb = 16'hfffe;
#10;
address_ina = 82;
address_inb = 83;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 84;
address_inb = 85;
data_ina = 16'h1;
data_inb = 16'h2;
#10;
address_ina = 86;
address_inb = 87;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 88;
address_inb = 89;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 90;
address_inb = 91;
data_ina = 16'h1;
data_inb = 16'h2;
#10;
address_ina = 92;
address_inb = 93;
data_ina = 16'h1;
data_inb = 16'hfffe;
#10;
address_ina = 94;
address_inb = 95;
data_ina = 16'h0;
data_inb = 16'hfffe;
#10;
address_ina = 96;
address_inb = 97;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 98;
address_inb = 99;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 100;
address_inb = 101;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 102;
address_inb = 103;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 104;
address_inb = 105;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 106;
address_inb = 107;
data_ina = 16'hfffe;
data_inb = 16'h2;
#10;
address_ina = 108;
address_inb = 109;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 110;
address_inb = 111;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 112;
address_inb = 113;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 114;
address_inb = 115;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 116;
address_inb = 117;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 118;
address_inb = 119;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 120;
address_inb = 121;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 122;
address_inb = 123;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 124;
address_inb = 125;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 126;
address_inb = 127;
data_ina = 16'h2;
data_inb = 16'hfffd;
#10;
address_ina = 128;
address_inb = 129;
data_ina = 16'h1;
data_inb = 16'h3;
#10;
address_ina = 130;
address_inb = 131;
data_ina = 16'h1;
data_inb = 16'h2;
#10;
address_ina = 132;
address_inb = 133;
data_ina = 16'hfffd;
data_inb = 16'h0;
#10;
address_ina = 134;
address_inb = 135;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 136;
address_inb = 137;
data_ina = 16'hfffd;
data_inb = 16'h0;
#10;
address_ina = 138;
address_inb = 139;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 140;
address_inb = 141;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 142;
address_inb = 143;
data_ina = 16'h2;
data_inb = 16'h1;
#10;
address_ina = 144;
address_inb = 145;
data_ina = 16'hfffe;
data_inb = 16'h0;
#10;
address_ina = 146;
address_inb = 147;
data_ina = 16'h1;
data_inb = 16'hfffe;
#10;
address_ina = 148;
address_inb = 149;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 150;
address_inb = 151;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 152;
address_inb = 153;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 154;
address_inb = 155;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 156;
address_inb = 157;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 158;
address_inb = 159;
data_ina = 16'h2;
data_inb = 16'hffff;
#10;
address_ina = 160;
address_inb = 161;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 162;
address_inb = 163;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 164;
address_inb = 165;
data_ina = 16'hffff;
data_inb = 16'hfffe;
#10;
address_ina = 166;
address_inb = 167;
data_ina = 16'h2;
data_inb = 16'hfffe;
#10;
address_ina = 168;
address_inb = 169;
data_ina = 16'h0;
data_inb = 16'h3;
#10;
address_ina = 170;
address_inb = 171;
data_ina = 16'h3;
data_inb = 16'hfffd;
#10;
address_ina = 172;
address_inb = 173;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 174;
address_inb = 175;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 176;
address_inb = 177;
data_ina = 16'h2;
data_inb = 16'h3;
#10;
address_ina = 178;
address_inb = 179;
data_ina = 16'h1;
data_inb = 16'h2;
#10;
address_ina = 180;
address_inb = 181;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 182;
address_inb = 183;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 184;
address_inb = 185;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 186;
address_inb = 187;
data_ina = 16'h1;
data_inb = 16'h2;
#10;
address_ina = 188;
address_inb = 189;
data_ina = 16'h2;
data_inb = 16'h1;
#10;
address_ina = 190;
address_inb = 191;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 192;
address_inb = 193;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 194;
address_inb = 195;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 196;
address_inb = 197;
data_ina = 16'h2;
data_inb = 16'hffff;
#10;
address_ina = 198;
address_inb = 199;
data_ina = 16'h0;
data_inb = 16'hfffe;
#10;
address_ina = 200;
address_inb = 201;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 202;
address_inb = 203;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 204;
address_inb = 205;
data_ina = 16'hfffe;
data_inb = 16'hfffe;
#10;
address_ina = 206;
address_inb = 207;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 208;
address_inb = 209;
data_ina = 16'hfffe;
data_inb = 16'h1;
#10;
address_ina = 210;
address_inb = 211;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 212;
address_inb = 213;
data_ina = 16'h1;
data_inb = 16'hfffe;
#10;
address_ina = 214;
address_inb = 215;
data_ina = 16'hffff;
data_inb = 16'hfffe;
#10;
address_ina = 216;
address_inb = 217;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 218;
address_inb = 219;
data_ina = 16'h0;
data_inb = 16'hfffe;
#10;
address_ina = 220;
address_inb = 221;
data_ina = 16'h2;
data_inb = 16'h3;
#10;
address_ina = 222;
address_inb = 223;
data_ina = 16'h0;
data_inb = 16'h2;
#10;
address_ina = 224;
address_inb = 225;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 226;
address_inb = 227;
data_ina = 16'hfffe;
data_inb = 16'hffff;
#10;
address_ina = 228;
address_inb = 229;
data_ina = 16'hfffd;
data_inb = 16'h0;
#10;
address_ina = 230;
address_inb = 231;
data_ina = 16'hfffe;
data_inb = 16'h2;
#10;
address_ina = 232;
address_inb = 233;
data_ina = 16'h3;
data_inb = 16'h0;
#10;
address_ina = 234;
address_inb = 235;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 236;
address_inb = 237;
data_ina = 16'hffff;
data_inb = 16'h2;
#10;
address_ina = 238;
address_inb = 239;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 240;
address_inb = 241;
data_ina = 16'h2;
data_inb = 16'h0;
#10;
address_ina = 242;
address_inb = 243;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 244;
address_inb = 245;
data_ina = 16'h2;
data_inb = 16'hffff;
#10;
address_ina = 246;
address_inb = 247;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 248;
address_inb = 249;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 250;
address_inb = 251;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 252;
address_inb = 253;
data_ina = 16'h2;
data_inb = 16'h0;
#10;
address_ina = 254;
address_inb = 255;
data_ina = 16'h0;
data_inb = 16'h3;
#10;
        wait(init_done);
        #30
        we = 0;
        // Start processing
         
		  #38000

        start = 0;



//        wait (wr_req);
//		  wait (!wr_req);
//		   rd_req = 1;
		  wait(done);
		  #20000
rd_req = 1;
        #70 
		  start = 1;
		 #80 
wait(rd_empty)
rd_req = 0;

$display("Finished the NTT test Number %d",test_num);
////Begin test number #5//////////////
rst = 1;

//#1000
start = 1;
mode = 0; //NTT 0 // INTT 1

// Reset for a few clock cycles

#1000

rst = 0;
test_num = test_num + 1;
#1000
we = 1;
address_ina = 0;
address_inb = 1;
data_ina = 16'h2;
data_inb = 16'h1;
#10;
address_ina = 2;
address_inb = 3;
data_ina = 16'hfffe;
data_inb = 16'hffff;
#10;
address_ina = 4;
address_inb = 5;
data_ina = 16'h2;
data_inb = 16'h1;
#10;
address_ina = 6;
address_inb = 7;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 8;
address_inb = 9;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 10;
address_inb = 11;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 12;
address_inb = 13;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 14;
address_inb = 15;
data_ina = 16'h1;
data_inb = 16'hfffe;
#10;
address_ina = 16;
address_inb = 17;
data_ina = 16'h2;
data_inb = 16'hfffe;
#10;
address_ina = 18;
address_inb = 19;
data_ina = 16'hfffe;
data_inb = 16'h1;
#10;
address_ina = 20;
address_inb = 21;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 22;
address_inb = 23;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 24;
address_inb = 25;
data_ina = 16'h0;
data_inb = 16'hfffe;
#10;
address_ina = 26;
address_inb = 27;
data_ina = 16'h2;
data_inb = 16'hffff;
#10;
address_ina = 28;
address_inb = 29;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 30;
address_inb = 31;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 32;
address_inb = 33;
data_ina = 16'h2;
data_inb = 16'hffff;
#10;
address_ina = 34;
address_inb = 35;
data_ina = 16'h2;
data_inb = 16'h1;
#10;
address_ina = 36;
address_inb = 37;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 38;
address_inb = 39;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 40;
address_inb = 41;
data_ina = 16'hfffe;
data_inb = 16'h0;
#10;
address_ina = 42;
address_inb = 43;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 44;
address_inb = 45;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 46;
address_inb = 47;
data_ina = 16'hfffe;
data_inb = 16'h1;
#10;
address_ina = 48;
address_inb = 49;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 50;
address_inb = 51;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 52;
address_inb = 53;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 54;
address_inb = 55;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 56;
address_inb = 57;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 58;
address_inb = 59;
data_ina = 16'h2;
data_inb = 16'h0;
#10;
address_ina = 60;
address_inb = 61;
data_ina = 16'h2;
data_inb = 16'h0;
#10;
address_ina = 62;
address_inb = 63;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 64;
address_inb = 65;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 66;
address_inb = 67;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 68;
address_inb = 69;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 70;
address_inb = 71;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 72;
address_inb = 73;
data_ina = 16'hfffe;
data_inb = 16'h1;
#10;
address_ina = 74;
address_inb = 75;
data_ina = 16'hfffd;
data_inb = 16'hffff;
#10;
address_ina = 76;
address_inb = 77;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 78;
address_inb = 79;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 80;
address_inb = 81;
data_ina = 16'h3;
data_inb = 16'h1;
#10;
address_ina = 82;
address_inb = 83;
data_ina = 16'h0;
data_inb = 16'h2;
#10;
address_ina = 84;
address_inb = 85;
data_ina = 16'h1;
data_inb = 16'h2;
#10;
address_ina = 86;
address_inb = 87;
data_ina = 16'hfffe;
data_inb = 16'h1;
#10;
address_ina = 88;
address_inb = 89;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 90;
address_inb = 91;
data_ina = 16'hfffe;
data_inb = 16'hffff;
#10;
address_ina = 92;
address_inb = 93;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 94;
address_inb = 95;
data_ina = 16'h0;
data_inb = 16'hfffe;
#10;
address_ina = 96;
address_inb = 97;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 98;
address_inb = 99;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 100;
address_inb = 101;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 102;
address_inb = 103;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 104;
address_inb = 105;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 106;
address_inb = 107;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 108;
address_inb = 109;
data_ina = 16'hfffd;
data_inb = 16'h0;
#10;
address_ina = 110;
address_inb = 111;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 112;
address_inb = 113;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 114;
address_inb = 115;
data_ina = 16'h1;
data_inb = 16'hfffe;
#10;
address_ina = 116;
address_inb = 117;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 118;
address_inb = 119;
data_ina = 16'hfffe;
data_inb = 16'hffff;
#10;
address_ina = 120;
address_inb = 121;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 122;
address_inb = 123;
data_ina = 16'hfffe;
data_inb = 16'h0;
#10;
address_ina = 124;
address_inb = 125;
data_ina = 16'h2;
data_inb = 16'h0;
#10;
address_ina = 126;
address_inb = 127;
data_ina = 16'h0;
data_inb = 16'hfffe;
#10;
address_ina = 128;
address_inb = 129;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 130;
address_inb = 131;
data_ina = 16'hfffe;
data_inb = 16'hffff;
#10;
address_ina = 132;
address_inb = 133;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 134;
address_inb = 135;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 136;
address_inb = 137;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 138;
address_inb = 139;
data_ina = 16'h1;
data_inb = 16'hfffd;
#10;
address_ina = 140;
address_inb = 141;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 142;
address_inb = 143;
data_ina = 16'h2;
data_inb = 16'h1;
#10;
address_ina = 144;
address_inb = 145;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 146;
address_inb = 147;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 148;
address_inb = 149;
data_ina = 16'h0;
data_inb = 16'hfffe;
#10;
address_ina = 150;
address_inb = 151;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 152;
address_inb = 153;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 154;
address_inb = 155;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 156;
address_inb = 157;
data_ina = 16'h0;
data_inb = 16'hfffe;
#10;
address_ina = 158;
address_inb = 159;
data_ina = 16'hffff;
data_inb = 16'hfffe;
#10;
address_ina = 160;
address_inb = 161;
data_ina = 16'h0;
data_inb = 16'h2;
#10;
address_ina = 162;
address_inb = 163;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 164;
address_inb = 165;
data_ina = 16'h2;
data_inb = 16'hfffd;
#10;
address_ina = 166;
address_inb = 167;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 168;
address_inb = 169;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 170;
address_inb = 171;
data_ina = 16'hfffe;
data_inb = 16'h1;
#10;
address_ina = 172;
address_inb = 173;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 174;
address_inb = 175;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 176;
address_inb = 177;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 178;
address_inb = 179;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 180;
address_inb = 181;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 182;
address_inb = 183;
data_ina = 16'hffff;
data_inb = 16'hfffe;
#10;
address_ina = 184;
address_inb = 185;
data_ina = 16'h0;
data_inb = 16'hfffe;
#10;
address_ina = 186;
address_inb = 187;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 188;
address_inb = 189;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 190;
address_inb = 191;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 192;
address_inb = 193;
data_ina = 16'h2;
data_inb = 16'h1;
#10;
address_ina = 194;
address_inb = 195;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 196;
address_inb = 197;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 198;
address_inb = 199;
data_ina = 16'hfffe;
data_inb = 16'h1;
#10;
address_ina = 200;
address_inb = 201;
data_ina = 16'hffff;
data_inb = 16'hfffe;
#10;
address_ina = 202;
address_inb = 203;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 204;
address_inb = 205;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 206;
address_inb = 207;
data_ina = 16'hfffe;
data_inb = 16'hffff;
#10;
address_ina = 208;
address_inb = 209;
data_ina = 16'hfffe;
data_inb = 16'h0;
#10;
address_ina = 210;
address_inb = 211;
data_ina = 16'hfffe;
data_inb = 16'hfffe;
#10;
address_ina = 212;
address_inb = 213;
data_ina = 16'hfffe;
data_inb = 16'h1;
#10;
address_ina = 214;
address_inb = 215;
data_ina = 16'h2;
data_inb = 16'h1;
#10;
address_ina = 216;
address_inb = 217;
data_ina = 16'h2;
data_inb = 16'hffff;
#10;
address_ina = 218;
address_inb = 219;
data_ina = 16'hffff;
data_inb = 16'hfffe;
#10;
address_ina = 220;
address_inb = 221;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 222;
address_inb = 223;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 224;
address_inb = 225;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 226;
address_inb = 227;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 228;
address_inb = 229;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 230;
address_inb = 231;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 232;
address_inb = 233;
data_ina = 16'h0;
data_inb = 16'h2;
#10;
address_ina = 234;
address_inb = 235;
data_ina = 16'h0;
data_inb = 16'h3;
#10;
address_ina = 236;
address_inb = 237;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 238;
address_inb = 239;
data_ina = 16'h1;
data_inb = 16'hfffe;
#10;
address_ina = 240;
address_inb = 241;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 242;
address_inb = 243;
data_ina = 16'hfffe;
data_inb = 16'hffff;
#10;
address_ina = 244;
address_inb = 245;
data_ina = 16'h0;
data_inb = 16'h2;
#10;
address_ina = 246;
address_inb = 247;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 248;
address_inb = 249;
data_ina = 16'hffff;
data_inb = 16'h3;
#10;
address_ina = 250;
address_inb = 251;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 252;
address_inb = 253;
data_ina = 16'h0;
data_inb = 16'hfffe;
#10;
address_ina = 254;
address_inb = 255;
data_ina = 16'h3;
data_inb = 16'h1;
#10;
        wait(init_done);
        #30
        we = 0;
        // Start processing
         
		  #38000

        start = 0;



//        wait (wr_req);
//		  wait (!wr_req);
//		   rd_req = 1;
		  wait(done);
		  #20000
rd_req = 1;
        #70 
		  start = 1;
		 #80 
wait(rd_empty)
rd_req = 0;

$display("Finished the NTT test Number %d",test_num);
////Begin test number #6//////////////
rst = 1;

//#1000
start = 1;
mode = 1; //NTT 0 // INTT 1

// Reset for a few clock cycles

#1000

rst = 0;
test_num = test_num + 1;
#1000
we = 1;
address_ina = 0;
address_inb = 1;
data_ina = 16'h410;
data_inb = 16'hf9e2;
#10;
address_ina = 2;
address_inb = 3;
data_ina = 16'h3be;
data_inb = 16'h43e;
#10;
address_ina = 4;
address_inb = 5;
data_ina = 16'h321;
data_inb = 16'h3f2;
#10;
address_ina = 6;
address_inb = 7;
data_ina = 16'hfac5;
data_inb = 16'h255;
#10;
address_ina = 8;
address_inb = 9;
data_ina = 16'hfe2b;
data_inb = 16'hff3d;
#10;
address_ina = 10;
address_inb = 11;
data_ina = 16'h420;
data_inb = 16'hfec1;
#10;
address_ina = 12;
address_inb = 13;
data_ina = 16'h215;
data_inb = 16'hfebe;
#10;
address_ina = 14;
address_inb = 15;
data_ina = 16'hfa07;
data_inb = 16'hfb98;
#10;
address_ina = 16;
address_inb = 17;
data_ina = 16'hff9a;
data_inb = 16'h41c;
#10;
address_ina = 18;
address_inb = 19;
data_ina = 16'hfcc0;
data_inb = 16'h17;
#10;
address_ina = 20;
address_inb = 21;
data_ina = 16'hfab0;
data_inb = 16'h2d8;
#10;
address_ina = 22;
address_inb = 23;
data_ina = 16'h2e3;
data_inb = 16'h665;
#10;
address_ina = 24;
address_inb = 25;
data_ina = 16'hfd2b;
data_inb = 16'h394;
#10;
address_ina = 26;
address_inb = 27;
data_ina = 16'hf98e;
data_inb = 16'h23c;
#10;
address_ina = 28;
address_inb = 29;
data_ina = 16'h560;
data_inb = 16'h313;
#10;
address_ina = 30;
address_inb = 31;
data_ina = 16'h203;
data_inb = 16'hfcd1;
#10;
address_ina = 32;
address_inb = 33;
data_ina = 16'h634;
data_inb = 16'hffcc;
#10;
address_ina = 34;
address_inb = 35;
data_ina = 16'hfeb6;
data_inb = 16'hfcc7;
#10;
address_ina = 36;
address_inb = 37;
data_ina = 16'hfa06;
data_inb = 16'hf98d;
#10;
address_ina = 38;
address_inb = 39;
data_ina = 16'h5fe;
data_inb = 16'hfcc4;
#10;
address_ina = 40;
address_inb = 41;
data_ina = 16'hfec6;
data_inb = 16'hfadd;
#10;
address_ina = 42;
address_inb = 43;
data_ina = 16'h92;
data_inb = 16'h25e;
#10;
address_ina = 44;
address_inb = 45;
data_ina = 16'h203;
data_inb = 16'hfbea;
#10;
address_ina = 46;
address_inb = 47;
data_ina = 16'h1b7;
data_inb = 16'hfc35;
#10;
address_ina = 48;
address_inb = 49;
data_ina = 16'h2db;
data_inb = 16'h156;
#10;
address_ina = 50;
address_inb = 51;
data_ina = 16'h4d5;
data_inb = 16'h40;
#10;
address_ina = 52;
address_inb = 53;
data_ina = 16'h1b;
data_inb = 16'hff7a;
#10;
address_ina = 54;
address_inb = 55;
data_ina = 16'h366;
data_inb = 16'hfa55;
#10;
address_ina = 56;
address_inb = 57;
data_ina = 16'h29c;
data_inb = 16'hfd96;
#10;
address_ina = 58;
address_inb = 59;
data_ina = 16'h515;
data_inb = 16'hfcd3;
#10;
address_ina = 60;
address_inb = 61;
data_ina = 16'h341;
data_inb = 16'h3ed;
#10;
address_ina = 62;
address_inb = 63;
data_ina = 16'h2e5;
data_inb = 16'h5a2;
#10;
address_ina = 64;
address_inb = 65;
data_ina = 16'h1e0;
data_inb = 16'hf9e3;
#10;
address_ina = 66;
address_inb = 67;
data_ina = 16'hfd01;
data_inb = 16'h262;
#10;
address_ina = 68;
address_inb = 69;
data_ina = 16'h42d;
data_inb = 16'hffed;
#10;
address_ina = 70;
address_inb = 71;
data_ina = 16'hfa45;
data_inb = 16'h2dd;
#10;
address_ina = 72;
address_inb = 73;
data_ina = 16'hffac;
data_inb = 16'h2a;
#10;
address_ina = 74;
address_inb = 75;
data_ina = 16'hfd4d;
data_inb = 16'h5a8;
#10;
address_ina = 76;
address_inb = 77;
data_ina = 16'hfd9c;
data_inb = 16'hff36;
#10;
address_ina = 78;
address_inb = 79;
data_ina = 16'h158;
data_inb = 16'hfbf3;
#10;
address_ina = 80;
address_inb = 81;
data_ina = 16'h676;
data_inb = 16'hfb11;
#10;
address_ina = 82;
address_inb = 83;
data_ina = 16'hfbd0;
data_inb = 16'h235;
#10;
address_ina = 84;
address_inb = 85;
data_ina = 16'h354;
data_inb = 16'h74;
#10;
address_ina = 86;
address_inb = 87;
data_ina = 16'hfdf7;
data_inb = 16'hfa56;
#10;
address_ina = 88;
address_inb = 89;
data_ina = 16'hfc60;
data_inb = 16'hfa5d;
#10;
address_ina = 90;
address_inb = 91;
data_ina = 16'hfddd;
data_inb = 16'h37f;
#10;
address_ina = 92;
address_inb = 93;
data_ina = 16'hff80;
data_inb = 16'hfba5;
#10;
address_ina = 94;
address_inb = 95;
data_ina = 16'h4c3;
data_inb = 16'hfa4c;
#10;
address_ina = 96;
address_inb = 97;
data_ina = 16'h51b;
data_inb = 16'hfe6d;
#10;
address_ina = 98;
address_inb = 99;
data_ina = 16'h53f;
data_inb = 16'hfe1c;
#10;
address_ina = 100;
address_inb = 101;
data_ina = 16'h1a0;
data_inb = 16'hf9fb;
#10;
address_ina = 102;
address_inb = 103;
data_ina = 16'h5b;
data_inb = 16'hfdb7;
#10;
address_ina = 104;
address_inb = 105;
data_ina = 16'ha3;
data_inb = 16'h3bc;
#10;
address_ina = 106;
address_inb = 107;
data_ina = 16'hfe2b;
data_inb = 16'hf9a5;
#10;
address_ina = 108;
address_inb = 109;
data_ina = 16'hfa79;
data_inb = 16'h4cd;
#10;
address_ina = 110;
address_inb = 111;
data_ina = 16'hfaac;
data_inb = 16'hfce2;
#10;
address_ina = 112;
address_inb = 113;
data_ina = 16'hfabb;
data_inb = 16'hfa83;
#10;
address_ina = 114;
address_inb = 115;
data_ina = 16'h124;
data_inb = 16'hfb1b;
#10;
address_ina = 116;
address_inb = 117;
data_ina = 16'hfe3d;
data_inb = 16'h65d;
#10;
address_ina = 118;
address_inb = 119;
data_ina = 16'h15d;
data_inb = 16'hff55;
#10;
address_ina = 120;
address_inb = 121;
data_ina = 16'h1ac;
data_inb = 16'hf4;
#10;
address_ina = 122;
address_inb = 123;
data_ina = 16'hfac2;
data_inb = 16'hee;
#10;
address_ina = 124;
address_inb = 125;
data_ina = 16'hfd7c;
data_inb = 16'h528;
#10;
address_ina = 126;
address_inb = 127;
data_ina = 16'hbc;
data_inb = 16'h17c;
#10;
address_ina = 128;
address_inb = 129;
data_ina = 16'h5e6;
data_inb = 16'hfb05;
#10;
address_ina = 130;
address_inb = 131;
data_ina = 16'h481;
data_inb = 16'h232;
#10;
address_ina = 132;
address_inb = 133;
data_ina = 16'hfc80;
data_inb = 16'hfdd3;
#10;
address_ina = 134;
address_inb = 135;
data_ina = 16'h6a;
data_inb = 16'h21f;
#10;
address_ina = 136;
address_inb = 137;
data_ina = 16'h5e5;
data_inb = 16'h1ff;
#10;
address_ina = 138;
address_inb = 139;
data_ina = 16'h377;
data_inb = 16'hfc81;
#10;
address_ina = 140;
address_inb = 141;
data_ina = 16'hfabe;
data_inb = 16'hfd73;
#10;
address_ina = 142;
address_inb = 143;
data_ina = 16'h5e;
data_inb = 16'he7;
#10;
address_ina = 144;
address_inb = 145;
data_ina = 16'h562;
data_inb = 16'h8;
#10;
address_ina = 146;
address_inb = 147;
data_ina = 16'h40a;
data_inb = 16'h9c;
#10;
address_ina = 148;
address_inb = 149;
data_ina = 16'h7;
data_inb = 16'h5ef;
#10;
address_ina = 150;
address_inb = 151;
data_ina = 16'hfbdd;
data_inb = 16'hfb00;
#10;
address_ina = 152;
address_inb = 153;
data_ina = 16'hfd29;
data_inb = 16'hfa94;
#10;
address_ina = 154;
address_inb = 155;
data_ina = 16'h134;
data_inb = 16'hfe63;
#10;
address_ina = 156;
address_inb = 157;
data_ina = 16'hfeb0;
data_inb = 16'h401;
#10;
address_ina = 158;
address_inb = 159;
data_ina = 16'hfb33;
data_inb = 16'hf9be;
#10;
address_ina = 160;
address_inb = 161;
data_ina = 16'h2fc;
data_inb = 16'hffdd;
#10;
address_ina = 162;
address_inb = 163;
data_ina = 16'hfb4d;
data_inb = 16'hfaf5;
#10;
address_ina = 164;
address_inb = 165;
data_ina = 16'h11e;
data_inb = 16'h1c5;
#10;
address_ina = 166;
address_inb = 167;
data_ina = 16'hfae6;
data_inb = 16'hc6;
#10;
address_ina = 168;
address_inb = 169;
data_ina = 16'hfd4e;
data_inb = 16'hfae6;
#10;
address_ina = 170;
address_inb = 171;
data_ina = 16'h35f;
data_inb = 16'h25b;
#10;
address_ina = 172;
address_inb = 173;
data_ina = 16'h2db;
data_inb = 16'h10c;
#10;
address_ina = 174;
address_inb = 175;
data_ina = 16'hfb6c;
data_inb = 16'hfa91;
#10;
address_ina = 176;
address_inb = 177;
data_ina = 16'h17d;
data_inb = 16'hfbbd;
#10;
address_ina = 178;
address_inb = 179;
data_ina = 16'h8c;
data_inb = 16'hff60;
#10;
address_ina = 180;
address_inb = 181;
data_ina = 16'hf9ea;
data_inb = 16'h620;
#10;
address_ina = 182;
address_inb = 183;
data_ina = 16'h1d1;
data_inb = 16'h22c;
#10;
address_ina = 184;
address_inb = 185;
data_ina = 16'h2a7;
data_inb = 16'h66;
#10;
address_ina = 186;
address_inb = 187;
data_ina = 16'hffd2;
data_inb = 16'hfc6b;
#10;
address_ina = 188;
address_inb = 189;
data_ina = 16'hff84;
data_inb = 16'hfcec;
#10;
address_ina = 190;
address_inb = 191;
data_ina = 16'h447;
data_inb = 16'hfa93;
#10;
address_ina = 192;
address_inb = 193;
data_ina = 16'h412;
data_inb = 16'hfae7;
#10;
address_ina = 194;
address_inb = 195;
data_ina = 16'hfb10;
data_inb = 16'hfc21;
#10;
address_ina = 196;
address_inb = 197;
data_ina = 16'h323;
data_inb = 16'h649;
#10;
address_ina = 198;
address_inb = 199;
data_ina = 16'hfee4;
data_inb = 16'hfeb5;
#10;
address_ina = 200;
address_inb = 201;
data_ina = 16'h441;
data_inb = 16'h21a;
#10;
address_ina = 202;
address_inb = 203;
data_ina = 16'h395;
data_inb = 16'heb;
#10;
address_ina = 204;
address_inb = 205;
data_ina = 16'hfca3;
data_inb = 16'h2f0;
#10;
address_ina = 206;
address_inb = 207;
data_ina = 16'h593;
data_inb = 16'hfa36;
#10;
address_ina = 208;
address_inb = 209;
data_ina = 16'hfac5;
data_inb = 16'hff18;
#10;
address_ina = 210;
address_inb = 211;
data_ina = 16'h288;
data_inb = 16'hfe04;
#10;
address_ina = 212;
address_inb = 213;
data_ina = 16'hfb92;
data_inb = 16'hfe33;
#10;
address_ina = 214;
address_inb = 215;
data_ina = 16'hfaad;
data_inb = 16'hfb26;
#10;
address_ina = 216;
address_inb = 217;
data_ina = 16'hff11;
data_inb = 16'hfb40;
#10;
address_ina = 218;
address_inb = 219;
data_ina = 16'h38;
data_inb = 16'hfa68;
#10;
address_ina = 220;
address_inb = 221;
data_ina = 16'hfd12;
data_inb = 16'hfa27;
#10;
address_ina = 222;
address_inb = 223;
data_ina = 16'h4e1;
data_inb = 16'h3e5;
#10;
address_ina = 224;
address_inb = 225;
data_ina = 16'hf990;
data_inb = 16'h317;
#10;
address_ina = 226;
address_inb = 227;
data_ina = 16'hf98e;
data_inb = 16'h53f;
#10;
address_ina = 228;
address_inb = 229;
data_ina = 16'hfa55;
data_inb = 16'h524;
#10;
address_ina = 230;
address_inb = 231;
data_ina = 16'hfd77;
data_inb = 16'h7;
#10;
address_ina = 232;
address_inb = 233;
data_ina = 16'hfe84;
data_inb = 16'h212;
#10;
address_ina = 234;
address_inb = 235;
data_ina = 16'hfbe2;
data_inb = 16'hfd33;
#10;
address_ina = 236;
address_inb = 237;
data_ina = 16'hfde4;
data_inb = 16'h98;
#10;
address_ina = 238;
address_inb = 239;
data_ina = 16'hfc36;
data_inb = 16'hfd85;
#10;
address_ina = 240;
address_inb = 241;
data_ina = 16'h325;
data_inb = 16'h37a;
#10;
address_ina = 242;
address_inb = 243;
data_ina = 16'hfa98;
data_inb = 16'hfbcb;
#10;
address_ina = 244;
address_inb = 245;
data_ina = 16'h12c;
data_inb = 16'h33f;
#10;
address_ina = 246;
address_inb = 247;
data_ina = 16'hfcde;
data_inb = 16'h407;
#10;
address_ina = 248;
address_inb = 249;
data_ina = 16'h520;
data_inb = 16'hfb70;
#10;
address_ina = 250;
address_inb = 251;
data_ina = 16'hff95;
data_inb = 16'h5e6;
#10;
address_ina = 252;
address_inb = 253;
data_ina = 16'hff84;
data_inb = 16'h166;
#10;
address_ina = 254;
address_inb = 255;
data_ina = 16'h66b;
data_inb = 16'h477;
#10;
        wait(init_done);
        #30
        we = 0;
        // Start processing
         
		  #38000

        start = 0;



//        wait (wr_req);
//		  wait (!wr_req);
//		   rd_req = 1;
		  wait(done);
		  #20000
rd_req = 1;
        #70 
		  start = 1;
		 #80 
wait(rd_empty)
rd_req = 0;

$display("Finished the NTT test Number %d",test_num);
////Begin test number #7//////////////
rst = 1;

//#1000
start = 1;
mode = 1; //NTT 0 // INTT 1

// Reset for a few clock cycles

#1000

rst = 0;
test_num = test_num + 1;
#1000
we = 1;
address_ina = 0;
address_inb = 1;
data_ina = 16'hfe35;
data_inb = 16'h378;
#10;
address_ina = 2;
address_inb = 3;
data_ina = 16'h455;
data_inb = 16'hfed6;
#10;
address_ina = 4;
address_inb = 5;
data_ina = 16'h62e;
data_inb = 16'hfaec;
#10;
address_ina = 6;
address_inb = 7;
data_ina = 16'hfe8d;
data_inb = 16'hfe7f;
#10;
address_ina = 8;
address_inb = 9;
data_ina = 16'hfe97;
data_inb = 16'hfbac;
#10;
address_ina = 10;
address_inb = 11;
data_ina = 16'hf9eb;
data_inb = 16'h65a;
#10;
address_ina = 12;
address_inb = 13;
data_ina = 16'hfd5b;
data_inb = 16'h57;
#10;
address_ina = 14;
address_inb = 15;
data_ina = 16'h460;
data_inb = 16'hf9ae;
#10;
address_ina = 16;
address_inb = 17;
data_ina = 16'h217;
data_inb = 16'h28a;
#10;
address_ina = 18;
address_inb = 19;
data_ina = 16'h436;
data_inb = 16'h36d;
#10;
address_ina = 20;
address_inb = 21;
data_ina = 16'h594;
data_inb = 16'h5d6;
#10;
address_ina = 22;
address_inb = 23;
data_ina = 16'hff50;
data_inb = 16'h1e0;
#10;
address_ina = 24;
address_inb = 25;
data_ina = 16'hfe0a;
data_inb = 16'hfdc3;
#10;
address_ina = 26;
address_inb = 27;
data_ina = 16'hfe7a;
data_inb = 16'hf9f3;
#10;
address_ina = 28;
address_inb = 29;
data_ina = 16'hfa10;
data_inb = 16'hf9b3;
#10;
address_ina = 30;
address_inb = 31;
data_ina = 16'hfa4a;
data_inb = 16'h2b8;
#10;
address_ina = 32;
address_inb = 33;
data_ina = 16'hff93;
data_inb = 16'hfe15;
#10;
address_ina = 34;
address_inb = 35;
data_ina = 16'h271;
data_inb = 16'hf9bf;
#10;
address_ina = 36;
address_inb = 37;
data_ina = 16'h579;
data_inb = 16'hff02;
#10;
address_ina = 38;
address_inb = 39;
data_ina = 16'h47e;
data_inb = 16'hfaed;
#10;
address_ina = 40;
address_inb = 41;
data_ina = 16'h548;
data_inb = 16'h427;
#10;
address_ina = 42;
address_inb = 43;
data_ina = 16'h1ac;
data_inb = 16'h608;
#10;
address_ina = 44;
address_inb = 45;
data_ina = 16'h6b;
data_inb = 16'hfcdb;
#10;
address_ina = 46;
address_inb = 47;
data_ina = 16'h1e6;
data_inb = 16'hfd4e;
#10;
address_ina = 48;
address_inb = 49;
data_ina = 16'hfe36;
data_inb = 16'hbd;
#10;
address_ina = 50;
address_inb = 51;
data_ina = 16'h42e;
data_inb = 16'h36f;
#10;
address_ina = 52;
address_inb = 53;
data_ina = 16'h3ca;
data_inb = 16'h1;
#10;
address_ina = 54;
address_inb = 55;
data_ina = 16'h473;
data_inb = 16'h5ce;
#10;
address_ina = 56;
address_inb = 57;
data_ina = 16'h79;
data_inb = 16'hf9e7;
#10;
address_ina = 58;
address_inb = 59;
data_ina = 16'hfb1d;
data_inb = 16'hff51;
#10;
address_ina = 60;
address_inb = 61;
data_ina = 16'h32c;
data_inb = 16'h4fc;
#10;
address_ina = 62;
address_inb = 63;
data_ina = 16'h8f;
data_inb = 16'hfe55;
#10;
address_ina = 64;
address_inb = 65;
data_ina = 16'h13f;
data_inb = 16'hfbe0;
#10;
address_ina = 66;
address_inb = 67;
data_ina = 16'hfc37;
data_inb = 16'h223;
#10;
address_ina = 68;
address_inb = 69;
data_ina = 16'h149;
data_inb = 16'hf2;
#10;
address_ina = 70;
address_inb = 71;
data_ina = 16'hfef9;
data_inb = 16'h2d9;
#10;
address_ina = 72;
address_inb = 73;
data_ina = 16'hfa7f;
data_inb = 16'hfc55;
#10;
address_ina = 74;
address_inb = 75;
data_ina = 16'h2c;
data_inb = 16'hfbdd;
#10;
address_ina = 76;
address_inb = 77;
data_ina = 16'hffcf;
data_inb = 16'h2b2;
#10;
address_ina = 78;
address_inb = 79;
data_ina = 16'hfdd1;
data_inb = 16'h36;
#10;
address_ina = 80;
address_inb = 81;
data_ina = 16'h27d;
data_inb = 16'hfffe;
#10;
address_ina = 82;
address_inb = 83;
data_ina = 16'h5f5;
data_inb = 16'h43b;
#10;
address_ina = 84;
address_inb = 85;
data_ina = 16'hf994;
data_inb = 16'hfa55;
#10;
address_ina = 86;
address_inb = 87;
data_ina = 16'hfd6b;
data_inb = 16'hfe50;
#10;
address_ina = 88;
address_inb = 89;
data_ina = 16'h58d;
data_inb = 16'h44f;
#10;
address_ina = 90;
address_inb = 91;
data_ina = 16'h1ad;
data_inb = 16'hfd8f;
#10;
address_ina = 92;
address_inb = 93;
data_ina = 16'hffab;
data_inb = 16'hfa0e;
#10;
address_ina = 94;
address_inb = 95;
data_ina = 16'hff5b;
data_inb = 16'h17c;
#10;
address_ina = 96;
address_inb = 97;
data_ina = 16'hfb0b;
data_inb = 16'h622;
#10;
address_ina = 98;
address_inb = 99;
data_ina = 16'hfcdc;
data_inb = 16'h1df;
#10;
address_ina = 100;
address_inb = 101;
data_ina = 16'h2e5;
data_inb = 16'hf9be;
#10;
address_ina = 102;
address_inb = 103;
data_ina = 16'h3f;
data_inb = 16'hfbb2;
#10;
address_ina = 104;
address_inb = 105;
data_ina = 16'h3ef;
data_inb = 16'h1a4;
#10;
address_ina = 106;
address_inb = 107;
data_ina = 16'hfdb6;
data_inb = 16'h4e2;
#10;
address_ina = 108;
address_inb = 109;
data_ina = 16'hfbc3;
data_inb = 16'hfbc4;
#10;
address_ina = 110;
address_inb = 111;
data_ina = 16'hfef6;
data_inb = 16'hf9ee;
#10;
address_ina = 112;
address_inb = 113;
data_ina = 16'hf9d9;
data_inb = 16'hff25;
#10;
address_ina = 114;
address_inb = 115;
data_ina = 16'hf9c1;
data_inb = 16'h275;
#10;
address_ina = 116;
address_inb = 117;
data_ina = 16'h65f;
data_inb = 16'hfa25;
#10;
address_ina = 118;
address_inb = 119;
data_ina = 16'h549;
data_inb = 16'h124;
#10;
address_ina = 120;
address_inb = 121;
data_ina = 16'h285;
data_inb = 16'h430;
#10;
address_ina = 122;
address_inb = 123;
data_ina = 16'hfebd;
data_inb = 16'hfb24;
#10;
address_ina = 124;
address_inb = 125;
data_ina = 16'hfa3a;
data_inb = 16'hfb03;
#10;
address_ina = 126;
address_inb = 127;
data_ina = 16'hfef2;
data_inb = 16'hff2c;
#10;
address_ina = 128;
address_inb = 129;
data_ina = 16'h175;
data_inb = 16'hfc8d;
#10;
address_ina = 130;
address_inb = 131;
data_ina = 16'hf7;
data_inb = 16'hfc0c;
#10;
address_ina = 132;
address_inb = 133;
data_ina = 16'hfdfb;
data_inb = 16'h49a;
#10;
address_ina = 134;
address_inb = 135;
data_ina = 16'hfffb;
data_inb = 16'h5ac;
#10;
address_ina = 136;
address_inb = 137;
data_ina = 16'hfe8a;
data_inb = 16'hff37;
#10;
address_ina = 138;
address_inb = 139;
data_ina = 16'hfd7b;
data_inb = 16'hfe98;
#10;
address_ina = 140;
address_inb = 141;
data_ina = 16'h451;
data_inb = 16'h19a;
#10;
address_ina = 142;
address_inb = 143;
data_ina = 16'h5ae;
data_inb = 16'hfdef;
#10;
address_ina = 144;
address_inb = 145;
data_ina = 16'h495;
data_inb = 16'h55;
#10;
address_ina = 146;
address_inb = 147;
data_ina = 16'hfc74;
data_inb = 16'hfb6a;
#10;
address_ina = 148;
address_inb = 149;
data_ina = 16'hfa0d;
data_inb = 16'h40d;
#10;
address_ina = 150;
address_inb = 151;
data_ina = 16'hffe6;
data_inb = 16'h51e;
#10;
address_ina = 152;
address_inb = 153;
data_ina = 16'hfd17;
data_inb = 16'hff28;
#10;
address_ina = 154;
address_inb = 155;
data_ina = 16'hfd08;
data_inb = 16'hfac1;
#10;
address_ina = 156;
address_inb = 157;
data_ina = 16'hfb44;
data_inb = 16'hfe08;
#10;
address_ina = 158;
address_inb = 159;
data_ina = 16'h57;
data_inb = 16'hfae6;
#10;
address_ina = 160;
address_inb = 161;
data_ina = 16'hfb04;
data_inb = 16'hfdb8;
#10;
address_ina = 162;
address_inb = 163;
data_ina = 16'hfe58;
data_inb = 16'h2ba;
#10;
address_ina = 164;
address_inb = 165;
data_ina = 16'hfb75;
data_inb = 16'h4ed;
#10;
address_ina = 166;
address_inb = 167;
data_ina = 16'hff1c;
data_inb = 16'hfbba;
#10;
address_ina = 168;
address_inb = 169;
data_ina = 16'h55c;
data_inb = 16'h5cf;
#10;
address_ina = 170;
address_inb = 171;
data_ina = 16'hfd7d;
data_inb = 16'hfa08;
#10;
address_ina = 172;
address_inb = 173;
data_ina = 16'hfc5e;
data_inb = 16'h4c8;
#10;
address_ina = 174;
address_inb = 175;
data_ina = 16'h6a;
data_inb = 16'h2c;
#10;
address_ina = 176;
address_inb = 177;
data_ina = 16'hfc15;
data_inb = 16'h82;
#10;
address_ina = 178;
address_inb = 179;
data_ina = 16'hfaf8;
data_inb = 16'h3ef;
#10;
address_ina = 180;
address_inb = 181;
data_ina = 16'h30e;
data_inb = 16'h507;
#10;
address_ina = 182;
address_inb = 183;
data_ina = 16'h445;
data_inb = 16'hfc77;
#10;
address_ina = 184;
address_inb = 185;
data_ina = 16'hfdd5;
data_inb = 16'h353;
#10;
address_ina = 186;
address_inb = 187;
data_ina = 16'h53d;
data_inb = 16'hfdf4;
#10;
address_ina = 188;
address_inb = 189;
data_ina = 16'hfd55;
data_inb = 16'hfa3a;
#10;
address_ina = 190;
address_inb = 191;
data_ina = 16'h1b7;
data_inb = 16'hfcaf;
#10;
address_ina = 192;
address_inb = 193;
data_ina = 16'hfb55;
data_inb = 16'hfa4b;
#10;
address_ina = 194;
address_inb = 195;
data_ina = 16'hfbe6;
data_inb = 16'hfb12;
#10;
address_ina = 196;
address_inb = 197;
data_ina = 16'h82;
data_inb = 16'h654;
#10;
address_ina = 198;
address_inb = 199;
data_ina = 16'hff49;
data_inb = 16'hff48;
#10;
address_ina = 200;
address_inb = 201;
data_ina = 16'h158;
data_inb = 16'hfb15;
#10;
address_ina = 202;
address_inb = 203;
data_ina = 16'hfa01;
data_inb = 16'h2f4;
#10;
address_ina = 204;
address_inb = 205;
data_ina = 16'h4a5;
data_inb = 16'h3f0;
#10;
address_ina = 206;
address_inb = 207;
data_ina = 16'hfd82;
data_inb = 16'h582;
#10;
address_ina = 208;
address_inb = 209;
data_ina = 16'h28f;
data_inb = 16'h4be;
#10;
address_ina = 210;
address_inb = 211;
data_ina = 16'h223;
data_inb = 16'h5be;
#10;
address_ina = 212;
address_inb = 213;
data_ina = 16'h518;
data_inb = 16'h214;
#10;
address_ina = 214;
address_inb = 215;
data_ina = 16'hfa8e;
data_inb = 16'hfca1;
#10;
address_ina = 216;
address_inb = 217;
data_ina = 16'hfafd;
data_inb = 16'hff0b;
#10;
address_ina = 218;
address_inb = 219;
data_ina = 16'h2ec;
data_inb = 16'h443;
#10;
address_ina = 220;
address_inb = 221;
data_ina = 16'h264;
data_inb = 16'h504;
#10;
address_ina = 222;
address_inb = 223;
data_ina = 16'hfb77;
data_inb = 16'hfc75;
#10;
address_ina = 224;
address_inb = 225;
data_ina = 16'hfd1a;
data_inb = 16'hfff4;
#10;
address_ina = 226;
address_inb = 227;
data_ina = 16'hfc57;
data_inb = 16'hff63;
#10;
address_ina = 228;
address_inb = 229;
data_ina = 16'h422;
data_inb = 16'h61a;
#10;
address_ina = 230;
address_inb = 231;
data_ina = 16'hfb3d;
data_inb = 16'h2e8;
#10;
address_ina = 232;
address_inb = 233;
data_ina = 16'h5a3;
data_inb = 16'hfb7a;
#10;
address_ina = 234;
address_inb = 235;
data_ina = 16'hfae8;
data_inb = 16'h57;
#10;
address_ina = 236;
address_inb = 237;
data_ina = 16'hfde6;
data_inb = 16'hf9b4;
#10;
address_ina = 238;
address_inb = 239;
data_ina = 16'h15d;
data_inb = 16'h2d2;
#10;
address_ina = 240;
address_inb = 241;
data_ina = 16'h493;
data_inb = 16'h163;
#10;
address_ina = 242;
address_inb = 243;
data_ina = 16'h322;
data_inb = 16'hffe4;
#10;
address_ina = 244;
address_inb = 245;
data_ina = 16'h466;
data_inb = 16'h144;
#10;
address_ina = 246;
address_inb = 247;
data_ina = 16'h366;
data_inb = 16'h623;
#10;
address_ina = 248;
address_inb = 249;
data_ina = 16'h48b;
data_inb = 16'h482;
#10;
address_ina = 250;
address_inb = 251;
data_ina = 16'hfb56;
data_inb = 16'h4;
#10;
address_ina = 252;
address_inb = 253;
data_ina = 16'hfeef;
data_inb = 16'h216;
#10;
address_ina = 254;
address_inb = 255;
data_ina = 16'h168;
data_inb = 16'heb;
#10;
        wait(init_done);
        #30
        we = 0;
        // Start processing
         
		  #38000

        start = 0;



//        wait (wr_req);
//		  wait (!wr_req);
//		   rd_req = 1;
		  wait(done);
		  #20000
rd_req = 1;
        #70 
		  start = 1;
		 #80 
wait(rd_empty)
rd_req = 0;

$display("Finished the NTT test Number %d",test_num);
////Begin test number #8//////////////
rst = 1;

//#1000
start = 1;
mode = 1; //NTT 0 // INTT 1

// Reset for a few clock cycles

#1000

rst = 0;
test_num = test_num + 1;
#1000
we = 1;
address_ina = 0;
address_inb = 1;
data_ina = 16'hfd21;
data_inb = 16'h277;
#10;
address_ina = 2;
address_inb = 3;
data_ina = 16'h2e1;
data_inb = 16'hfb1f;
#10;
address_ina = 4;
address_inb = 5;
data_ina = 16'h5c6;
data_inb = 16'h132;
#10;
address_ina = 6;
address_inb = 7;
data_ina = 16'h4e2;
data_inb = 16'hc1;
#10;
address_ina = 8;
address_inb = 9;
data_ina = 16'hf9cb;
data_inb = 16'hfaf0;
#10;
address_ina = 10;
address_inb = 11;
data_ina = 16'hfef0;
data_inb = 16'hff0c;
#10;
address_ina = 12;
address_inb = 13;
data_ina = 16'h60;
data_inb = 16'h59;
#10;
address_ina = 14;
address_inb = 15;
data_ina = 16'hfa33;
data_inb = 16'h67b;
#10;
address_ina = 16;
address_inb = 17;
data_ina = 16'hfb8b;
data_inb = 16'hfd38;
#10;
address_ina = 18;
address_inb = 19;
data_ina = 16'hfa82;
data_inb = 16'hff;
#10;
address_ina = 20;
address_inb = 21;
data_ina = 16'h603;
data_inb = 16'h3fa;
#10;
address_ina = 22;
address_inb = 23;
data_ina = 16'hf999;
data_inb = 16'hfc01;
#10;
address_ina = 24;
address_inb = 25;
data_ina = 16'h2f2;
data_inb = 16'h159;
#10;
address_ina = 26;
address_inb = 27;
data_ina = 16'hfd0b;
data_inb = 16'h339;
#10;
address_ina = 28;
address_inb = 29;
data_ina = 16'hfa9e;
data_inb = 16'h505;
#10;
address_ina = 30;
address_inb = 31;
data_ina = 16'hfe7e;
data_inb = 16'hfdcc;
#10;
address_ina = 32;
address_inb = 33;
data_ina = 16'h34a;
data_inb = 16'hfb3f;
#10;
address_ina = 34;
address_inb = 35;
data_ina = 16'hfb6a;
data_inb = 16'h17a;
#10;
address_ina = 36;
address_inb = 37;
data_ina = 16'h33c;
data_inb = 16'h608;
#10;
address_ina = 38;
address_inb = 39;
data_ina = 16'h181;
data_inb = 16'hff88;
#10;
address_ina = 40;
address_inb = 41;
data_ina = 16'hfd7e;
data_inb = 16'hff1e;
#10;
address_ina = 42;
address_inb = 43;
data_ina = 16'h5be;
data_inb = 16'h580;
#10;
address_ina = 44;
address_inb = 45;
data_ina = 16'h66c;
data_inb = 16'hfaed;
#10;
address_ina = 46;
address_inb = 47;
data_ina = 16'h4a1;
data_inb = 16'hfd15;
#10;
address_ina = 48;
address_inb = 49;
data_ina = 16'hfff1;
data_inb = 16'hfb55;
#10;
address_ina = 50;
address_inb = 51;
data_ina = 16'h174;
data_inb = 16'hfc83;
#10;
address_ina = 52;
address_inb = 53;
data_ina = 16'hfe72;
data_inb = 16'hffa9;
#10;
address_ina = 54;
address_inb = 55;
data_ina = 16'hfdab;
data_inb = 16'h5b5;
#10;
address_ina = 56;
address_inb = 57;
data_ina = 16'hfcdd;
data_inb = 16'h1a8;
#10;
address_ina = 58;
address_inb = 59;
data_ina = 16'hfef2;
data_inb = 16'hfd41;
#10;
address_ina = 60;
address_inb = 61;
data_ina = 16'hfd75;
data_inb = 16'hfd52;
#10;
address_ina = 62;
address_inb = 63;
data_ina = 16'hfa16;
data_inb = 16'hfaee;
#10;
address_ina = 64;
address_inb = 65;
data_ina = 16'hff47;
data_inb = 16'h331;
#10;
address_ina = 66;
address_inb = 67;
data_ina = 16'hfe8c;
data_inb = 16'hfea3;
#10;
address_ina = 68;
address_inb = 69;
data_ina = 16'hffa3;
data_inb = 16'hba;
#10;
address_ina = 70;
address_inb = 71;
data_ina = 16'h19;
data_inb = 16'hfad0;
#10;
address_ina = 72;
address_inb = 73;
data_ina = 16'hff5c;
data_inb = 16'h4e4;
#10;
address_ina = 74;
address_inb = 75;
data_ina = 16'h2e;
data_inb = 16'h645;
#10;
address_ina = 76;
address_inb = 77;
data_ina = 16'hfebf;
data_inb = 16'hffaa;
#10;
address_ina = 78;
address_inb = 79;
data_ina = 16'hfee0;
data_inb = 16'h42;
#10;
address_ina = 80;
address_inb = 81;
data_ina = 16'h361;
data_inb = 16'hffec;
#10;
address_ina = 82;
address_inb = 83;
data_ina = 16'hff68;
data_inb = 16'hfb49;
#10;
address_ina = 84;
address_inb = 85;
data_ina = 16'hfa28;
data_inb = 16'h20;
#10;
address_ina = 86;
address_inb = 87;
data_ina = 16'hfdd1;
data_inb = 16'hfc77;
#10;
address_ina = 88;
address_inb = 89;
data_ina = 16'hfdd5;
data_inb = 16'hfd40;
#10;
address_ina = 90;
address_inb = 91;
data_ina = 16'hfa94;
data_inb = 16'hfaab;
#10;
address_ina = 92;
address_inb = 93;
data_ina = 16'hf9a1;
data_inb = 16'hff9c;
#10;
address_ina = 94;
address_inb = 95;
data_ina = 16'h2f9;
data_inb = 16'hfc77;
#10;
address_ina = 96;
address_inb = 97;
data_ina = 16'hfc13;
data_inb = 16'h442;
#10;
address_ina = 98;
address_inb = 99;
data_ina = 16'hfbc9;
data_inb = 16'hfbcf;
#10;
address_ina = 100;
address_inb = 101;
data_ina = 16'h13f;
data_inb = 16'hfc34;
#10;
address_ina = 102;
address_inb = 103;
data_ina = 16'h1ed;
data_inb = 16'h104;
#10;
address_ina = 104;
address_inb = 105;
data_ina = 16'h1c2;
data_inb = 16'hfad7;
#10;
address_ina = 106;
address_inb = 107;
data_ina = 16'hfbb2;
data_inb = 16'hfc38;
#10;
address_ina = 108;
address_inb = 109;
data_ina = 16'hfe33;
data_inb = 16'hfb40;
#10;
address_ina = 110;
address_inb = 111;
data_ina = 16'hfaba;
data_inb = 16'h12;
#10;
address_ina = 112;
address_inb = 113;
data_ina = 16'hf98b;
data_inb = 16'h44c;
#10;
address_ina = 114;
address_inb = 115;
data_ina = 16'h310;
data_inb = 16'hff4e;
#10;
address_ina = 116;
address_inb = 117;
data_ina = 16'hfb5a;
data_inb = 16'h32e;
#10;
address_ina = 118;
address_inb = 119;
data_ina = 16'hfb6f;
data_inb = 16'hfbf1;
#10;
address_ina = 120;
address_inb = 121;
data_ina = 16'hff4c;
data_inb = 16'hfe0d;
#10;
address_ina = 122;
address_inb = 123;
data_ina = 16'hfe0a;
data_inb = 16'hfdd3;
#10;
address_ina = 124;
address_inb = 125;
data_ina = 16'hfaaa;
data_inb = 16'hfe15;
#10;
address_ina = 126;
address_inb = 127;
data_ina = 16'h412;
data_inb = 16'hfc2f;
#10;
address_ina = 128;
address_inb = 129;
data_ina = 16'hfa41;
data_inb = 16'hf9cd;
#10;
address_ina = 130;
address_inb = 131;
data_ina = 16'h32a;
data_inb = 16'h5e5;
#10;
address_ina = 132;
address_inb = 133;
data_ina = 16'h297;
data_inb = 16'h1a2;
#10;
address_ina = 134;
address_inb = 135;
data_ina = 16'hfb90;
data_inb = 16'h60f;
#10;
address_ina = 136;
address_inb = 137;
data_ina = 16'hfecb;
data_inb = 16'h27b;
#10;
address_ina = 138;
address_inb = 139;
data_ina = 16'hfaf2;
data_inb = 16'h310;
#10;
address_ina = 140;
address_inb = 141;
data_ina = 16'h390;
data_inb = 16'hfe6d;
#10;
address_ina = 142;
address_inb = 143;
data_ina = 16'h4cf;
data_inb = 16'h427;
#10;
address_ina = 144;
address_inb = 145;
data_ina = 16'hf9e2;
data_inb = 16'h134;
#10;
address_ina = 146;
address_inb = 147;
data_ina = 16'hfc28;
data_inb = 16'h565;
#10;
address_ina = 148;
address_inb = 149;
data_ina = 16'hfacd;
data_inb = 16'hfc70;
#10;
address_ina = 150;
address_inb = 151;
data_ina = 16'h3c2;
data_inb = 16'hfd7e;
#10;
address_ina = 152;
address_inb = 153;
data_ina = 16'hfd32;
data_inb = 16'hf9f7;
#10;
address_ina = 154;
address_inb = 155;
data_ina = 16'h560;
data_inb = 16'hf9ab;
#10;
address_ina = 156;
address_inb = 157;
data_ina = 16'hfabe;
data_inb = 16'h5b7;
#10;
address_ina = 158;
address_inb = 159;
data_ina = 16'hfd2b;
data_inb = 16'hfe93;
#10;
address_ina = 160;
address_inb = 161;
data_ina = 16'h49;
data_inb = 16'h2d3;
#10;
address_ina = 162;
address_inb = 163;
data_ina = 16'h51a;
data_inb = 16'h348;
#10;
address_ina = 164;
address_inb = 165;
data_ina = 16'h23f;
data_inb = 16'h3cb;
#10;
address_ina = 166;
address_inb = 167;
data_ina = 16'hfb27;
data_inb = 16'hff08;
#10;
address_ina = 168;
address_inb = 169;
data_ina = 16'hfb41;
data_inb = 16'hfd0e;
#10;
address_ina = 170;
address_inb = 171;
data_ina = 16'hff7f;
data_inb = 16'h661;
#10;
address_ina = 172;
address_inb = 173;
data_ina = 16'had;
data_inb = 16'h54;
#10;
address_ina = 174;
address_inb = 175;
data_ina = 16'hfffd;
data_inb = 16'hfb61;
#10;
address_ina = 176;
address_inb = 177;
data_ina = 16'hfd29;
data_inb = 16'hfabb;
#10;
address_ina = 178;
address_inb = 179;
data_ina = 16'hd8;
data_inb = 16'hfeff;
#10;
address_ina = 180;
address_inb = 181;
data_ina = 16'h445;
data_inb = 16'hfddb;
#10;
address_ina = 182;
address_inb = 183;
data_ina = 16'he3;
data_inb = 16'h520;
#10;
address_ina = 184;
address_inb = 185;
data_ina = 16'hfc35;
data_inb = 16'hff26;
#10;
address_ina = 186;
address_inb = 187;
data_ina = 16'hfab5;
data_inb = 16'h208;
#10;
address_ina = 188;
address_inb = 189;
data_ina = 16'hfe3d;
data_inb = 16'h191;
#10;
address_ina = 190;
address_inb = 191;
data_ina = 16'hfbb2;
data_inb = 16'hfab5;
#10;
address_ina = 192;
address_inb = 193;
data_ina = 16'hfa85;
data_inb = 16'h494;
#10;
address_ina = 194;
address_inb = 195;
data_ina = 16'hfb7a;
data_inb = 16'h463;
#10;
address_ina = 196;
address_inb = 197;
data_ina = 16'hfb6b;
data_inb = 16'h101;
#10;
address_ina = 198;
address_inb = 199;
data_ina = 16'h15d;
data_inb = 16'h593;
#10;
address_ina = 200;
address_inb = 201;
data_ina = 16'h29e;
data_inb = 16'hfa67;
#10;
address_ina = 202;
address_inb = 203;
data_ina = 16'h25d;
data_inb = 16'hfd87;
#10;
address_ina = 204;
address_inb = 205;
data_ina = 16'hef;
data_inb = 16'h373;
#10;
address_ina = 206;
address_inb = 207;
data_ina = 16'h210;
data_inb = 16'h5da;
#10;
address_ina = 208;
address_inb = 209;
data_ina = 16'hfd8b;
data_inb = 16'hff8d;
#10;
address_ina = 210;
address_inb = 211;
data_ina = 16'hf985;
data_inb = 16'hfa38;
#10;
address_ina = 212;
address_inb = 213;
data_ina = 16'h1e4;
data_inb = 16'h65a;
#10;
address_ina = 214;
address_inb = 215;
data_ina = 16'hfa19;
data_inb = 16'h23d;
#10;
address_ina = 216;
address_inb = 217;
data_ina = 16'h249;
data_inb = 16'hfcd4;
#10;
address_ina = 218;
address_inb = 219;
data_ina = 16'hfc8d;
data_inb = 16'hfa0f;
#10;
address_ina = 220;
address_inb = 221;
data_ina = 16'h537;
data_inb = 16'hfa46;
#10;
address_ina = 222;
address_inb = 223;
data_ina = 16'hfd49;
data_inb = 16'hfecb;
#10;
address_ina = 224;
address_inb = 225;
data_ina = 16'h5c2;
data_inb = 16'hfe4a;
#10;
address_ina = 226;
address_inb = 227;
data_ina = 16'h174;
data_inb = 16'hfb0e;
#10;
address_ina = 228;
address_inb = 229;
data_ina = 16'h410;
data_inb = 16'hfe16;
#10;
address_ina = 230;
address_inb = 231;
data_ina = 16'h0;
data_inb = 16'h478;
#10;
address_ina = 232;
address_inb = 233;
data_ina = 16'h1bc;
data_inb = 16'h57d;
#10;
address_ina = 234;
address_inb = 235;
data_ina = 16'h3cc;
data_inb = 16'h275;
#10;
address_ina = 236;
address_inb = 237;
data_ina = 16'hfd2d;
data_inb = 16'hfd60;
#10;
address_ina = 238;
address_inb = 239;
data_ina = 16'h1dc;
data_inb = 16'h36c;
#10;
address_ina = 240;
address_inb = 241;
data_ina = 16'hfac3;
data_inb = 16'h132;
#10;
address_ina = 242;
address_inb = 243;
data_ina = 16'h568;
data_inb = 16'h67;
#10;
address_ina = 244;
address_inb = 245;
data_ina = 16'h3de;
data_inb = 16'hfc10;
#10;
address_ina = 246;
address_inb = 247;
data_ina = 16'h156;
data_inb = 16'h4a5;
#10;
address_ina = 248;
address_inb = 249;
data_ina = 16'hfe84;
data_inb = 16'h5c1;
#10;
address_ina = 250;
address_inb = 251;
data_ina = 16'hfab5;
data_inb = 16'h53d;
#10;
address_ina = 252;
address_inb = 253;
data_ina = 16'hfc4b;
data_inb = 16'hfd07;
#10;
address_ina = 254;
address_inb = 255;
data_ina = 16'hfb6a;
data_inb = 16'h15d;
#10;
        wait(init_done);
        #30
        we = 0;
        // Start processing
         
		  #38000

        start = 0;



//        wait (wr_req);
//		  wait (!wr_req);
//		   rd_req = 1;
		  wait(done);
		  #20000
rd_req = 1;
        #70 
		  start = 1;
		 #80 
wait(rd_empty)
rd_req = 0;

$display("Finished the NTT test Number %d",test_num);
////Begin test number #9//////////////
rst = 1;

//#1000
start = 1;
mode = 0; //NTT 0 // INTT 1

// Reset for a few clock cycles

#1000

rst = 0;
test_num = test_num + 1;
#1000
we = 1;
address_ina = 0;
address_inb = 1;
data_ina = 16'h8b9;
data_inb = 16'h7cf;
#10;
address_ina = 2;
address_inb = 3;
data_ina = 16'h21f;
data_inb = 16'h989;
#10;
address_ina = 4;
address_inb = 5;
data_ina = 16'ha9;
data_inb = 16'h2ab;
#10;
address_ina = 6;
address_inb = 7;
data_ina = 16'h754;
data_inb = 16'ha49;
#10;
address_ina = 8;
address_inb = 9;
data_ina = 16'hced;
data_inb = 16'h538;
#10;
address_ina = 10;
address_inb = 11;
data_ina = 16'h6ef;
data_inb = 16'h781;
#10;
address_ina = 12;
address_inb = 13;
data_ina = 16'h6dc;
data_inb = 16'h911;
#10;
address_ina = 14;
address_inb = 15;
data_ina = 16'h31c;
data_inb = 16'h246;
#10;
address_ina = 16;
address_inb = 17;
data_ina = 16'hc78;
data_inb = 16'h8e4;
#10;
address_ina = 18;
address_inb = 19;
data_ina = 16'hced;
data_inb = 16'h88f;
#10;
address_ina = 20;
address_inb = 21;
data_ina = 16'haf2;
data_inb = 16'h344;
#10;
address_ina = 22;
address_inb = 23;
data_ina = 16'h892;
data_inb = 16'h36b;
#10;
address_ina = 24;
address_inb = 25;
data_ina = 16'haff;
data_inb = 16'h58;
#10;
address_ina = 26;
address_inb = 27;
data_ina = 16'h8b3;
data_inb = 16'h1bd;
#10;
address_ina = 28;
address_inb = 29;
data_ina = 16'h72;
data_inb = 16'h589;
#10;
address_ina = 30;
address_inb = 31;
data_ina = 16'h114;
data_inb = 16'hca3;
#10;
address_ina = 32;
address_inb = 33;
data_ina = 16'h75;
data_inb = 16'h24c;
#10;
address_ina = 34;
address_inb = 35;
data_ina = 16'h632;
data_inb = 16'h744;
#10;
address_ina = 36;
address_inb = 37;
data_ina = 16'h80a;
data_inb = 16'h11b;
#10;
address_ina = 38;
address_inb = 39;
data_ina = 16'h569;
data_inb = 16'h60b;
#10;
address_ina = 40;
address_inb = 41;
data_ina = 16'haf2;
data_inb = 16'h7cf;
#10;
address_ina = 42;
address_inb = 43;
data_ina = 16'hc72;
data_inb = 16'h189;
#10;
address_ina = 44;
address_inb = 45;
data_ina = 16'hb57;
data_inb = 16'h38b;
#10;
address_ina = 46;
address_inb = 47;
data_ina = 16'h3c6;
data_inb = 16'h80d;
#10;
address_ina = 48;
address_inb = 49;
data_ina = 16'h3ac;
data_inb = 16'h76b;
#10;
address_ina = 50;
address_inb = 51;
data_ina = 16'h8b9;
data_inb = 16'h93f;
#10;
address_ina = 52;
address_inb = 53;
data_ina = 16'h5fe;
data_inb = 16'h10b;
#10;
address_ina = 54;
address_inb = 55;
data_ina = 16'h892;
data_inb = 16'h2ab;
#10;
address_ina = 56;
address_inb = 57;
data_ina = 16'hb4a;
data_inb = 16'h51b;
#10;
address_ina = 58;
address_inb = 59;
data_ina = 16'h36b;
data_inb = 16'h6dc;
#10;
address_ina = 60;
address_inb = 61;
data_ina = 16'h555;
data_inb = 16'h703;
#10;
address_ina = 62;
address_inb = 63;
data_ina = 16'h636;
data_inb = 16'h42e;
#10;
address_ina = 64;
address_inb = 65;
data_ina = 16'h6cf;
data_inb = 16'h53f;
#10;
address_ina = 66;
address_inb = 67;
data_ina = 16'hb19;
data_inb = 16'h3e3;
#10;
address_ina = 68;
address_inb = 69;
data_ina = 16'h48f;
data_inb = 16'hcf4;
#10;
address_ina = 70;
address_inb = 71;
data_ina = 16'h9c;
data_inb = 16'he7;
#10;
address_ina = 72;
address_inb = 73;
data_ina = 16'hc68;
data_inb = 16'h1c1;
#10;
address_ina = 74;
address_inb = 75;
data_ina = 16'h2be;
data_inb = 16'h996;
#10;
address_ina = 76;
address_inb = 77;
data_ina = 16'h632;
data_inb = 16'h615;
#10;
address_ina = 78;
address_inb = 79;
data_ina = 16'h8da;
data_inb = 16'h68;
#10;
address_ina = 80;
address_inb = 81;
data_ina = 16'h236;
data_inb = 16'h4a6;
#10;
address_ina = 82;
address_inb = 83;
data_ina = 16'h2e2;
data_inb = 16'hc37;
#10;
address_ina = 84;
address_inb = 85;
data_ina = 16'h69b;
data_inb = 16'h236;
#10;
address_ina = 86;
address_inb = 87;
data_ina = 16'h95f;
data_inb = 16'h77e;
#10;
address_ina = 88;
address_inb = 89;
data_ina = 16'h40a;
data_inb = 16'h33a;
#10;
address_ina = 90;
address_inb = 91;
data_ina = 16'h9c7;
data_inb = 16'h75a;
#10;
address_ina = 92;
address_inb = 93;
data_ina = 16'h407;
data_inb = 16'ha60;
#10;
address_ina = 94;
address_inb = 95;
data_ina = 16'ha08;
data_inb = 16'hc92;
#10;
address_ina = 96;
address_inb = 97;
data_ina = 16'hcd3;
data_inb = 16'h7ed;
#10;
address_ina = 98;
address_inb = 99;
data_ina = 16'h2db;
data_inb = 16'h489;
#10;
address_ina = 100;
address_inb = 101;
data_ina = 16'hac2;
data_inb = 16'h256;
#10;
address_ina = 102;
address_inb = 103;
data_ina = 16'hbb2;
data_inb = 16'h7c9;
#10;
address_ina = 104;
address_inb = 105;
data_ina = 16'h336;
data_inb = 16'h865;
#10;
address_ina = 106;
address_inb = 107;
data_ina = 16'hb10;
data_inb = 16'h9e8;
#10;
address_ina = 108;
address_inb = 109;
data_ina = 16'h5b7;
data_inb = 16'h7bc;
#10;
address_ina = 110;
address_inb = 111;
data_ina = 16'hc5b;
data_inb = 16'h4f4;
#10;
address_ina = 112;
address_inb = 113;
data_ina = 16'h78e;
data_inb = 16'h788;
#10;
address_ina = 114;
address_inb = 115;
data_ina = 16'hcb0;
data_inb = 16'h528;
#10;
address_ina = 116;
address_inb = 117;
data_ina = 16'hb19;
data_inb = 16'h5e4;
#10;
address_ina = 118;
address_inb = 119;
data_ina = 16'h9f;
data_inb = 16'hb13;
#10;
address_ina = 120;
address_inb = 121;
data_ina = 16'h7d3;
data_inb = 16'h507;
#10;
address_ina = 122;
address_inb = 123;
data_ina = 16'h5b0;
data_inb = 16'h59a;
#10;
address_ina = 124;
address_inb = 125;
data_ina = 16'he0;
data_inb = 16'h1eb;
#10;
address_ina = 126;
address_inb = 127;
data_ina = 16'hb23;
data_inb = 16'h2c8;
#10;
address_ina = 128;
address_inb = 129;
data_ina = 16'h5a0;
data_inb = 16'h525;
#10;
address_ina = 130;
address_inb = 131;
data_ina = 16'h24;
data_inb = 16'h521;
#10;
address_ina = 132;
address_inb = 133;
data_ina = 16'h670;
data_inb = 16'hcfa;
#10;
address_ina = 134;
address_inb = 135;
data_ina = 16'h7bf;
data_inb = 16'h125;
#10;
address_ina = 136;
address_inb = 137;
data_ina = 16'h42a;
data_inb = 16'h12e;
#10;
address_ina = 138;
address_inb = 139;
data_ina = 16'hd7;
data_inb = 16'hc9c;
#10;
address_ina = 140;
address_inb = 141;
data_ina = 16'h649;
data_inb = 16'h118;
#10;
address_ina = 142;
address_inb = 143;
data_ina = 16'h785;
data_inb = 16'h511;
#10;
address_ina = 144;
address_inb = 145;
data_ina = 16'h807;
data_inb = 16'h514;
#10;
address_ina = 146;
address_inb = 147;
data_ina = 16'h385;
data_inb = 16'h67a;
#10;
address_ina = 148;
address_inb = 149;
data_ina = 16'h407;
data_inb = 16'hb0;
#10;
address_ina = 150;
address_inb = 151;
data_ina = 16'h542;
data_inb = 16'h511;
#10;
address_ina = 152;
address_inb = 153;
data_ina = 16'hcf1;
data_inb = 16'hc34;
#10;
address_ina = 154;
address_inb = 155;
data_ina = 16'h125;
data_inb = 16'ha70;
#10;
address_ina = 156;
address_inb = 157;
data_ina = 16'ha02;
data_inb = 16'h737;
#10;
address_ina = 158;
address_inb = 159;
data_ina = 16'h263;
data_inb = 16'h30f;
#10;
address_ina = 160;
address_inb = 161;
data_ina = 16'h8dd;
data_inb = 16'h46b;
#10;
address_ina = 162;
address_inb = 163;
data_ina = 16'h6df;
data_inb = 16'h2e8;
#10;
address_ina = 164;
address_inb = 165;
data_ina = 16'hb81;
data_inb = 16'h990;
#10;
address_ina = 166;
address_inb = 167;
data_ina = 16'h684;
data_inb = 16'h562;
#10;
address_ina = 168;
address_inb = 169;
data_ina = 16'h767;
data_inb = 16'h6ae;
#10;
address_ina = 170;
address_inb = 171;
data_ina = 16'h21f;
data_inb = 16'h96c;
#10;
address_ina = 172;
address_inb = 173;
data_ina = 16'h190;
data_inb = 16'h455;
#10;
address_ina = 174;
address_inb = 175;
data_ina = 16'h12b;
data_inb = 16'h2d8;
#10;
address_ina = 176;
address_inb = 177;
data_ina = 16'hcb9;
data_inb = 16'h18d;
#10;
address_ina = 178;
address_inb = 179;
data_ina = 16'hc37;
data_inb = 16'hc6;
#10;
address_ina = 180;
address_inb = 181;
data_ina = 16'h6a1;
data_inb = 16'hcd;
#10;
address_ina = 182;
address_inb = 183;
data_ina = 16'hae2;
data_inb = 16'h407;
#10;
address_ina = 184;
address_inb = 185;
data_ina = 16'h344;
data_inb = 16'h1d1;
#10;
address_ina = 186;
address_inb = 187;
data_ina = 16'h132;
data_inb = 16'h882;
#10;
address_ina = 188;
address_inb = 189;
data_ina = 16'h7e0;
data_inb = 16'h771;
#10;
address_ina = 190;
address_inb = 191;
data_ina = 16'h361;
data_inb = 16'h142;
#10;
address_ina = 192;
address_inb = 193;
data_ina = 16'ha81;
data_inb = 16'hbd6;
#10;
address_ina = 194;
address_inb = 195;
data_ina = 16'h7f0;
data_inb = 16'had8;
#10;
address_ina = 196;
address_inb = 197;
data_ina = 16'h218;
data_inb = 16'h76b;
#10;
address_ina = 198;
address_inb = 199;
data_ina = 16'h9d8;
data_inb = 16'hb81;
#10;
address_ina = 200;
address_inb = 201;
data_ina = 16'h9b4;
data_inb = 16'h5b7;
#10;
address_ina = 202;
address_inb = 203;
data_ina = 16'h5fe;
data_inb = 16'h9eb;
#10;
address_ina = 204;
address_inb = 205;
data_ina = 16'h50b;
data_inb = 16'h392;
#10;
address_ina = 206;
address_inb = 207;
data_ina = 16'h330;
data_inb = 16'h807;
#10;
address_ina = 208;
address_inb = 209;
data_ina = 16'h986;
data_inb = 16'h6f9;
#10;
address_ina = 210;
address_inb = 211;
data_ina = 16'h7;
data_inb = 16'h236;
#10;
address_ina = 212;
address_inb = 213;
data_ina = 16'h6f9;
data_inb = 16'h468;
#10;
address_ina = 214;
address_inb = 215;
data_ina = 16'h632;
data_inb = 16'h336;
#10;
address_ina = 216;
address_inb = 217;
data_ina = 16'hbbf;
data_inb = 16'hc9c;
#10;
address_ina = 218;
address_inb = 219;
data_ina = 16'h37e;
data_inb = 16'h3fd;
#10;
address_ina = 220;
address_inb = 221;
data_ina = 16'h989;
data_inb = 16'h19a;
#10;
address_ina = 222;
address_inb = 223;
data_ina = 16'h7a2;
data_inb = 16'h91b;
#10;
address_ina = 224;
address_inb = 225;
data_ina = 16'habb;
data_inb = 16'hbc2;
#10;
address_ina = 226;
address_inb = 227;
data_ina = 16'h189;
data_inb = 16'h77e;
#10;
address_ina = 228;
address_inb = 229;
data_ina = 16'h7ed;
data_inb = 16'h263;
#10;
address_ina = 230;
address_inb = 231;
data_ina = 16'h2d2;
data_inb = 16'h2b4;
#10;
address_ina = 232;
address_inb = 233;
data_ina = 16'h21f;
data_inb = 16'h403;
#10;
address_ina = 234;
address_inb = 235;
data_ina = 16'h719;
data_inb = 16'h7a5;
#10;
address_ina = 236;
address_inb = 237;
data_ina = 16'h4fe;
data_inb = 16'h63c;
#10;
address_ina = 238;
address_inb = 239;
data_ina = 16'h20b;
data_inb = 16'he7;
#10;
address_ina = 240;
address_inb = 241;
data_ina = 16'hccd;
data_inb = 16'h280;
#10;
address_ina = 242;
address_inb = 243;
data_ina = 16'h1e8;
data_inb = 16'hcf7;
#10;
address_ina = 244;
address_inb = 245;
data_ina = 16'h60f;
data_inb = 16'h84b;
#10;
address_ina = 246;
address_inb = 247;
data_ina = 16'h9fb;
data_inb = 16'h605;
#10;
address_ina = 248;
address_inb = 249;
data_ina = 16'h9ff;
data_inb = 16'h643;
#10;
address_ina = 250;
address_inb = 251;
data_ina = 16'hbb5;
data_inb = 16'h878;
#10;
address_ina = 252;
address_inb = 253;
data_ina = 16'h193;
data_inb = 16'hca6;
#10;
address_ina = 254;
address_inb = 255;
data_ina = 16'h697;
data_inb = 16'h212;
#10;
        wait(init_done);
        #30
        we = 0;
        // Start processing
         
		  #38000

        start = 0;



//        wait (wr_req);
//		  wait (!wr_req);
//		   rd_req = 1;
		  wait(done);
		  #20000
rd_req = 1;
        #70 
		  start = 1;
		 #80 
wait(rd_empty)
rd_req = 0;

$display("Finished the NTT test Number %d",test_num);
////Begin test number #10//////////////
rst = 1;

//#1000
start = 1;
mode = 0; //NTT 0 // INTT 1

// Reset for a few clock cycles

#1000

rst = 0;
test_num = test_num + 1;
#1000
we = 1;
address_ina = 0;
address_inb = 1;
data_ina = 16'h834;
data_inb = 16'h4d0;
#10;
address_ina = 2;
address_inb = 3;
data_ina = 16'h5ad;
data_inb = 16'h559;
#10;
address_ina = 4;
address_inb = 5;
data_ina = 16'h3cc;
data_inb = 16'h193;
#10;
address_ina = 6;
address_inb = 7;
data_ina = 16'h72;
data_inb = 16'h4b9;
#10;
address_ina = 8;
address_inb = 9;
data_ina = 16'h7e3;
data_inb = 16'h25d;
#10;
address_ina = 10;
address_inb = 11;
data_ina = 16'hb6;
data_inb = 16'h36e;
#10;
address_ina = 12;
address_inb = 13;
data_ina = 16'h0;
data_inb = 16'h720;
#10;
address_ina = 14;
address_inb = 15;
data_ina = 16'hc92;
data_inb = 16'h13f;
#10;
address_ina = 16;
address_inb = 17;
data_ina = 16'h821;
data_inb = 16'h7dc;
#10;
address_ina = 18;
address_inb = 19;
data_ina = 16'h3c2;
data_inb = 16'hcac;
#10;
address_ina = 20;
address_inb = 21;
data_ina = 16'hc51;
data_inb = 16'h46f;
#10;
address_ina = 22;
address_inb = 23;
data_ina = 16'h694;
data_inb = 16'h7f3;
#10;
address_ina = 24;
address_inb = 25;
data_ina = 16'hcd0;
data_inb = 16'hb6b;
#10;
address_ina = 26;
address_inb = 27;
data_ina = 16'h3e9;
data_inb = 16'h4f7;
#10;
address_ina = 28;
address_inb = 29;
data_ina = 16'hbf3;
data_inb = 16'h5db;
#10;
address_ina = 30;
address_inb = 31;
data_ina = 16'hc5b;
data_inb = 16'ha36;
#10;
address_ina = 32;
address_inb = 33;
data_ina = 16'h444;
data_inb = 16'h3cc;
#10;
address_ina = 34;
address_inb = 35;
data_ina = 16'hc41;
data_inb = 16'hc9c;
#10;
address_ina = 36;
address_inb = 37;
data_ina = 16'h7f;
data_inb = 16'hcd3;
#10;
address_ina = 38;
address_inb = 39;
data_ina = 16'h650;
data_inb = 16'h8ea;
#10;
address_ina = 40;
address_inb = 41;
data_ina = 16'h771;
data_inb = 16'h35e;
#10;
address_ina = 42;
address_inb = 43;
data_ina = 16'h37b;
data_inb = 16'h8f1;
#10;
address_ina = 44;
address_inb = 45;
data_ina = 16'h458;
data_inb = 16'h6d2;
#10;
address_ina = 46;
address_inb = 47;
data_ina = 16'h9c1;
data_inb = 16'ha60;
#10;
address_ina = 48;
address_inb = 49;
data_ina = 16'hb9f;
data_inb = 16'h5f5;
#10;
address_ina = 50;
address_inb = 51;
data_ina = 16'h256;
data_inb = 16'h86b;
#10;
address_ina = 52;
address_inb = 53;
data_ina = 16'hb98;
data_inb = 16'h80a;
#10;
address_ina = 54;
address_inb = 55;
data_ina = 16'h132;
data_inb = 16'h79f;
#10;
address_ina = 56;
address_inb = 57;
data_ina = 16'hae9;
data_inb = 16'h851;
#10;
address_ina = 58;
address_inb = 59;
data_ina = 16'h180;
data_inb = 16'h37e;
#10;
address_ina = 60;
address_inb = 61;
data_ina = 16'h559;
data_inb = 16'h7f;
#10;
address_ina = 62;
address_inb = 63;
data_ina = 16'h2f9;
data_inb = 16'h785;
#10;
address_ina = 64;
address_inb = 65;
data_ina = 16'h751;
data_inb = 16'hcfa;
#10;
address_ina = 66;
address_inb = 67;
data_ina = 16'h681;
data_inb = 16'h99a;
#10;
address_ina = 68;
address_inb = 69;
data_ina = 16'h63f;
data_inb = 16'hb10;
#10;
address_ina = 70;
address_inb = 71;
data_ina = 16'h111;
data_inb = 16'h771;
#10;
address_ina = 72;
address_inb = 73;
data_ina = 16'h632;
data_inb = 16'h99;
#10;
address_ina = 74;
address_inb = 75;
data_ina = 16'h45b;
data_inb = 16'hcd3;
#10;
address_ina = 76;
address_inb = 77;
data_ina = 16'h650;
data_inb = 16'h1a;
#10;
address_ina = 78;
address_inb = 79;
data_ina = 16'hc37;
data_inb = 16'h62c;
#10;
address_ina = 80;
address_inb = 81;
data_ina = 16'h468;
data_inb = 16'h31c;
#10;
address_ina = 82;
address_inb = 83;
data_ina = 16'ha74;
data_inb = 16'h166;
#10;
address_ina = 84;
address_inb = 85;
data_ina = 16'ha8e;
data_inb = 16'h9cb;
#10;
address_ina = 86;
address_inb = 87;
data_ina = 16'h1d4;
data_inb = 16'h747;
#10;
address_ina = 88;
address_inb = 89;
data_ina = 16'ha36;
data_inb = 16'hc21;
#10;
address_ina = 90;
address_inb = 91;
data_ina = 16'h5ad;
data_inb = 16'h59a;
#10;
address_ina = 92;
address_inb = 93;
data_ina = 16'haa1;
data_inb = 16'h8a9;
#10;
address_ina = 94;
address_inb = 95;
data_ina = 16'h914;
data_inb = 16'hbcc;
#10;
address_ina = 96;
address_inb = 97;
data_ina = 16'h507;
data_inb = 16'h896;
#10;
address_ina = 98;
address_inb = 99;
data_ina = 16'h615;
data_inb = 16'h43b;
#10;
address_ina = 100;
address_inb = 101;
data_ina = 16'hccd;
data_inb = 16'hb0;
#10;
address_ina = 102;
address_inb = 103;
data_ina = 16'h4e0;
data_inb = 16'h5d1;
#10;
address_ina = 104;
address_inb = 105;
data_ina = 16'h85b;
data_inb = 16'haf9;
#10;
address_ina = 106;
address_inb = 107;
data_ina = 16'hacf;
data_inb = 16'h3bc;
#10;
address_ina = 108;
address_inb = 109;
data_ina = 16'hf7;
data_inb = 16'h656;
#10;
address_ina = 110;
address_inb = 111;
data_ina = 16'hce0;
data_inb = 16'h81d;
#10;
address_ina = 112;
address_inb = 113;
data_ina = 16'h142;
data_inb = 16'hb74;
#10;
address_ina = 114;
address_inb = 115;
data_ina = 16'hbf3;
data_inb = 16'h4ea;
#10;
address_ina = 116;
address_inb = 117;
data_ina = 16'h7e0;
data_inb = 16'h785;
#10;
address_ina = 118;
address_inb = 119;
data_ina = 16'h55;
data_inb = 16'h97c;
#10;
address_ina = 120;
address_inb = 121;
data_ina = 16'h44;
data_inb = 16'h6d2;
#10;
address_ina = 122;
address_inb = 123;
data_ina = 16'h69b;
data_inb = 16'hbf6;
#10;
address_ina = 124;
address_inb = 125;
data_ina = 16'hb7b;
data_inb = 16'h421;
#10;
address_ina = 126;
address_inb = 127;
data_ina = 16'h5e4;
data_inb = 16'ha9;
#10;
address_ina = 128;
address_inb = 129;
data_ina = 16'hbac;
data_inb = 16'h76e;
#10;
address_ina = 130;
address_inb = 131;
data_ina = 16'h865;
data_inb = 16'h788;
#10;
address_ina = 132;
address_inb = 133;
data_ina = 16'h5aa;
data_inb = 16'h6e2;
#10;
address_ina = 134;
address_inb = 135;
data_ina = 16'h496;
data_inb = 16'h28d;
#10;
address_ina = 136;
address_inb = 137;
data_ina = 16'hae2;
data_inb = 16'had5;
#10;
address_ina = 138;
address_inb = 139;
data_ina = 16'h81a;
data_inb = 16'h326;
#10;
address_ina = 140;
address_inb = 141;
data_ina = 16'h189;
data_inb = 16'h3cf;
#10;
address_ina = 142;
address_inb = 143;
data_ina = 16'h76b;
data_inb = 16'h277;
#10;
address_ina = 144;
address_inb = 145;
data_ina = 16'h9db;
data_inb = 16'h892;
#10;
address_ina = 146;
address_inb = 147;
data_ina = 16'hc6b;
data_inb = 16'h48;
#10;
address_ina = 148;
address_inb = 149;
data_ina = 16'h357;
data_inb = 16'ha56;
#10;
address_ina = 150;
address_inb = 151;
data_ina = 16'h28d;
data_inb = 16'h4e0;
#10;
address_ina = 152;
address_inb = 153;
data_ina = 16'had8;
data_inb = 16'h962;
#10;
address_ina = 154;
address_inb = 155;
data_ina = 16'h751;
data_inb = 16'hbb5;
#10;
address_ina = 156;
address_inb = 157;
data_ina = 16'hb16;
data_inb = 16'h85b;
#10;
address_ina = 158;
address_inb = 159;
data_ina = 16'h421;
data_inb = 16'h7a2;
#10;
address_ina = 160;
address_inb = 161;
data_ina = 16'h862;
data_inb = 16'hce7;
#10;
address_ina = 162;
address_inb = 163;
data_ina = 16'hc48;
data_inb = 16'hb9f;
#10;
address_ina = 164;
address_inb = 165;
data_ina = 16'h2c1;
data_inb = 16'ha0f;
#10;
address_ina = 166;
address_inb = 167;
data_ina = 16'h9f;
data_inb = 16'h990;
#10;
address_ina = 168;
address_inb = 169;
data_ina = 16'h966;
data_inb = 16'h518;
#10;
address_ina = 170;
address_inb = 171;
data_ina = 16'h50b;
data_inb = 16'h767;
#10;
address_ina = 172;
address_inb = 173;
data_ina = 16'hb20;
data_inb = 16'h5ca;
#10;
address_ina = 174;
address_inb = 175;
data_ina = 16'hbed;
data_inb = 16'h485;
#10;
address_ina = 176;
address_inb = 177;
data_ina = 16'hc0a;
data_inb = 16'h3b2;
#10;
address_ina = 178;
address_inb = 179;
data_ina = 16'h19a;
data_inb = 16'h179;
#10;
address_ina = 180;
address_inb = 181;
data_ina = 16'h78e;
data_inb = 16'h2bb;
#10;
address_ina = 182;
address_inb = 183;
data_ina = 16'h6ab;
data_inb = 16'h596;
#10;
address_ina = 184;
address_inb = 185;
data_ina = 16'h3f0;
data_inb = 16'h548;
#10;
address_ina = 186;
address_inb = 187;
data_ina = 16'hc2a;
data_inb = 16'h84e;
#10;
address_ina = 188;
address_inb = 189;
data_ina = 16'h3d3;
data_inb = 16'hc00;
#10;
address_ina = 190;
address_inb = 191;
data_ina = 16'h538;
data_inb = 16'h465;
#10;
address_ina = 192;
address_inb = 193;
data_ina = 16'h1b0;
data_inb = 16'h125;
#10;
address_ina = 194;
address_inb = 195;
data_ina = 16'h2d8;
data_inb = 16'h4cd;
#10;
address_ina = 196;
address_inb = 197;
data_ina = 16'hbd;
data_inb = 16'h3a8;
#10;
address_ina = 198;
address_inb = 199;
data_ina = 16'h253;
data_inb = 16'ha05;
#10;
address_ina = 200;
address_inb = 201;
data_ina = 16'h478;
data_inb = 16'h979;
#10;
address_ina = 202;
address_inb = 203;
data_ina = 16'hc17;
data_inb = 16'h12e;
#10;
address_ina = 204;
address_inb = 205;
data_ina = 16'h118;
data_inb = 16'h34;
#10;
address_ina = 206;
address_inb = 207;
data_ina = 16'hc21;
data_inb = 16'hc1d;
#10;
address_ina = 208;
address_inb = 209;
data_ina = 16'hc78;
data_inb = 16'h35e;
#10;
address_ina = 210;
address_inb = 211;
data_ina = 16'h99a;
data_inb = 16'h6dc;
#10;
address_ina = 212;
address_inb = 213;
data_ina = 16'h59d;
data_inb = 16'h4a9;
#10;
address_ina = 214;
address_inb = 215;
data_ina = 16'h643;
data_inb = 16'h3c6;
#10;
address_ina = 216;
address_inb = 217;
data_ina = 16'h518;
data_inb = 16'h309;
#10;
address_ina = 218;
address_inb = 219;
data_ina = 16'h90b;
data_inb = 16'h580;
#10;
address_ina = 220;
address_inb = 221;
data_ina = 16'haa4;
data_inb = 16'h54f;
#10;
address_ina = 222;
address_inb = 223;
data_ina = 16'haef;
data_inb = 16'h7a2;
#10;
address_ina = 224;
address_inb = 225;
data_ina = 16'h320;
data_inb = 16'hc10;
#10;
address_ina = 226;
address_inb = 227;
data_ina = 16'hc78;
data_inb = 16'h46b;
#10;
address_ina = 228;
address_inb = 229;
data_ina = 16'h37b;
data_inb = 16'h431;
#10;
address_ina = 230;
address_inb = 231;
data_ina = 16'h514;
data_inb = 16'h4fe;
#10;
address_ina = 232;
address_inb = 233;
data_ina = 16'hb09;
data_inb = 16'hbed;
#10;
address_ina = 234;
address_inb = 235;
data_ina = 16'hd0;
data_inb = 16'hac8;
#10;
address_ina = 236;
address_inb = 237;
data_ina = 16'h35a;
data_inb = 16'h9f8;
#10;
address_ina = 238;
address_inb = 239;
data_ina = 16'h608;
data_inb = 16'h82;
#10;
address_ina = 240;
address_inb = 241;
data_ina = 16'h788;
data_inb = 16'h48f;
#10;
address_ina = 242;
address_inb = 243;
data_ina = 16'h125;
data_inb = 16'h4c6;
#10;
address_ina = 244;
address_inb = 245;
data_ina = 16'h5de;
data_inb = 16'h697;
#10;
address_ina = 246;
address_inb = 247;
data_ina = 16'hcb6;
data_inb = 16'h367;
#10;
address_ina = 248;
address_inb = 249;
data_ina = 16'hb98;
data_inb = 16'h3d3;
#10;
address_ina = 250;
address_inb = 251;
data_ina = 16'h3e3;
data_inb = 16'h26d;
#10;
address_ina = 252;
address_inb = 253;
data_ina = 16'h205;
data_inb = 16'h5c7;
#10;
address_ina = 254;
address_inb = 255;
data_ina = 16'hac8;
data_inb = 16'h858;
#10;
        wait(init_done);
        #30
        we = 0;
        // Start processing
         
		  #38000

        start = 0;



//        wait (wr_req);
//		  wait (!wr_req);
//		   rd_req = 1;
		  wait(done);
		  #20000
rd_req = 1;
        #70 
		  start = 1;
		 #80 
wait(rd_empty)
rd_req = 0;

$display("Finished the NTT test Number %d",test_num);
////Begin test number #11//////////////
rst = 1;

//#1000
start = 1;
mode = 1; //NTT 0 // INTT 1

// Reset for a few clock cycles

#1000

rst = 0;
test_num = test_num + 1;
#1000
we = 1;
address_ina = 0;
address_inb = 1;
data_ina = 16'hfc86;
data_inb = 16'h3e0;
#10;
address_ina = 2;
address_inb = 3;
data_ina = 16'h3cd;
data_inb = 16'h93;
#10;
address_ina = 4;
address_inb = 5;
data_ina = 16'hfd8b;
data_inb = 16'h106;
#10;
address_ina = 6;
address_inb = 7;
data_ina = 16'h32a;
data_inb = 16'h6d;
#10;
address_ina = 8;
address_inb = 9;
data_ina = 16'h15;
data_inb = 16'hfa90;
#10;
address_ina = 10;
address_inb = 11;
data_ina = 16'hffe5;
data_inb = 16'hfca9;
#10;
address_ina = 12;
address_inb = 13;
data_ina = 16'h5da;
data_inb = 16'h209;
#10;
address_ina = 14;
address_inb = 15;
data_ina = 16'hfab4;
data_inb = 16'h1b;
#10;
address_ina = 16;
address_inb = 17;
data_ina = 16'h429;
data_inb = 16'hfb8a;
#10;
address_ina = 18;
address_inb = 19;
data_ina = 16'h641;
data_inb = 16'h548;
#10;
address_ina = 20;
address_inb = 21;
data_ina = 16'h2ab;
data_inb = 16'hfb14;
#10;
address_ina = 22;
address_inb = 23;
data_ina = 16'h60d;
data_inb = 16'h221;
#10;
address_ina = 24;
address_inb = 25;
data_ina = 16'hfa7e;
data_inb = 16'hfee7;
#10;
address_ina = 26;
address_inb = 27;
data_ina = 16'h3fb;
data_inb = 16'h455;
#10;
address_ina = 28;
address_inb = 29;
data_ina = 16'hff31;
data_inb = 16'h304;
#10;
address_ina = 30;
address_inb = 31;
data_ina = 16'h287;
data_inb = 16'hfeec;
#10;
address_ina = 32;
address_inb = 33;
data_ina = 16'hfb46;
data_inb = 16'h166;
#10;
address_ina = 34;
address_inb = 35;
data_ina = 16'h441;
data_inb = 16'hf980;
#10;
address_ina = 36;
address_inb = 37;
data_ina = 16'h5d7;
data_inb = 16'hff3e;
#10;
address_ina = 38;
address_inb = 39;
data_ina = 16'h426;
data_inb = 16'h5ca;
#10;
address_ina = 40;
address_inb = 41;
data_ina = 16'hfe9b;
data_inb = 16'hfaed;
#10;
address_ina = 42;
address_inb = 43;
data_ina = 16'h177;
data_inb = 16'h169;
#10;
address_ina = 44;
address_inb = 45;
data_ina = 16'h390;
data_inb = 16'hfae2;
#10;
address_ina = 46;
address_inb = 47;
data_ina = 16'h523;
data_inb = 16'hfad0;
#10;
address_ina = 48;
address_inb = 49;
data_ina = 16'h337;
data_inb = 16'h39b;
#10;
address_ina = 50;
address_inb = 51;
data_ina = 16'hf994;
data_inb = 16'h4c4;
#10;
address_ina = 52;
address_inb = 53;
data_ina = 16'hfbdd;
data_inb = 16'hfcd5;
#10;
address_ina = 54;
address_inb = 55;
data_ina = 16'hfc87;
data_inb = 16'h1d1;
#10;
address_ina = 56;
address_inb = 57;
data_ina = 16'hfaff;
data_inb = 16'hfbb2;
#10;
address_ina = 58;
address_inb = 59;
data_ina = 16'h68;
data_inb = 16'hfb60;
#10;
address_ina = 60;
address_inb = 61;
data_ina = 16'hc0;
data_inb = 16'h25;
#10;
address_ina = 62;
address_inb = 63;
data_ina = 16'hfae8;
data_inb = 16'h36f;
#10;
address_ina = 64;
address_inb = 65;
data_ina = 16'h8a;
data_inb = 16'h57a;
#10;
address_ina = 66;
address_inb = 67;
data_ina = 16'h588;
data_inb = 16'hfb60;
#10;
address_ina = 68;
address_inb = 69;
data_ina = 16'hfd94;
data_inb = 16'hfc57;
#10;
address_ina = 70;
address_inb = 71;
data_ina = 16'h192;
data_inb = 16'hfb60;
#10;
address_ina = 72;
address_inb = 73;
data_ina = 16'hfae6;
data_inb = 16'hfc5f;
#10;
address_ina = 74;
address_inb = 75;
data_ina = 16'hfc41;
data_inb = 16'h3b9;
#10;
address_ina = 76;
address_inb = 77;
data_ina = 16'h1eb;
data_inb = 16'hfeb6;
#10;
address_ina = 78;
address_inb = 79;
data_ina = 16'hfd67;
data_inb = 16'hfb8c;
#10;
address_ina = 80;
address_inb = 81;
data_ina = 16'hfd1f;
data_inb = 16'hfb41;
#10;
address_ina = 82;
address_inb = 83;
data_ina = 16'hfd47;
data_inb = 16'h593;
#10;
address_ina = 84;
address_inb = 85;
data_ina = 16'hfe7f;
data_inb = 16'hfc7f;
#10;
address_ina = 86;
address_inb = 87;
data_ina = 16'h407;
data_inb = 16'hfe86;
#10;
address_ina = 88;
address_inb = 89;
data_ina = 16'hfc9e;
data_inb = 16'h19d;
#10;
address_ina = 90;
address_inb = 91;
data_ina = 16'hfd23;
data_inb = 16'h4f7;
#10;
address_ina = 92;
address_inb = 93;
data_ina = 16'h5d4;
data_inb = 16'hfc69;
#10;
address_ina = 94;
address_inb = 95;
data_ina = 16'h134;
data_inb = 16'h5c6;
#10;
address_ina = 96;
address_inb = 97;
data_ina = 16'h494;
data_inb = 16'he;
#10;
address_ina = 98;
address_inb = 99;
data_ina = 16'hfca8;
data_inb = 16'h3fb;
#10;
address_ina = 100;
address_inb = 101;
data_ina = 16'h3a3;
data_inb = 16'hfbc1;
#10;
address_ina = 102;
address_inb = 103;
data_ina = 16'hfcaa;
data_inb = 16'hf9cf;
#10;
address_ina = 104;
address_inb = 105;
data_ina = 16'hfad6;
data_inb = 16'h390;
#10;
address_ina = 106;
address_inb = 107;
data_ina = 16'hfdee;
data_inb = 16'hbe;
#10;
address_ina = 108;
address_inb = 109;
data_ina = 16'hfb98;
data_inb = 16'hd8;
#10;
address_ina = 110;
address_inb = 111;
data_ina = 16'hffbb;
data_inb = 16'h490;
#10;
address_ina = 112;
address_inb = 113;
data_ina = 16'hffb5;
data_inb = 16'h41;
#10;
address_ina = 114;
address_inb = 115;
data_ina = 16'h321;
data_inb = 16'hfb36;
#10;
address_ina = 116;
address_inb = 117;
data_ina = 16'h191;
data_inb = 16'hfcd0;
#10;
address_ina = 118;
address_inb = 119;
data_ina = 16'hffd9;
data_inb = 16'hfc80;
#10;
address_ina = 120;
address_inb = 121;
data_ina = 16'he3;
data_inb = 16'hfbd7;
#10;
address_ina = 122;
address_inb = 123;
data_ina = 16'hfbae;
data_inb = 16'h5d0;
#10;
address_ina = 124;
address_inb = 125;
data_ina = 16'hfd79;
data_inb = 16'h386;
#10;
address_ina = 126;
address_inb = 127;
data_ina = 16'hfc7e;
data_inb = 16'hfe34;
#10;
address_ina = 128;
address_inb = 129;
data_ina = 16'h441;
data_inb = 16'hff60;
#10;
address_ina = 130;
address_inb = 131;
data_ina = 16'hc8;
data_inb = 16'h365;
#10;
address_ina = 132;
address_inb = 133;
data_ina = 16'h5bf;
data_inb = 16'h139;
#10;
address_ina = 134;
address_inb = 135;
data_ina = 16'hfce4;
data_inb = 16'hfefb;
#10;
address_ina = 136;
address_inb = 137;
data_ina = 16'h83;
data_inb = 16'hfd8f;
#10;
address_ina = 138;
address_inb = 139;
data_ina = 16'h4d4;
data_inb = 16'h8e;
#10;
address_ina = 140;
address_inb = 141;
data_ina = 16'h33c;
data_inb = 16'h27d;
#10;
address_ina = 142;
address_inb = 143;
data_ina = 16'hfe4c;
data_inb = 16'h595;
#10;
address_ina = 144;
address_inb = 145;
data_ina = 16'h265;
data_inb = 16'h490;
#10;
address_ina = 146;
address_inb = 147;
data_ina = 16'hfb55;
data_inb = 16'h3a;
#10;
address_ina = 148;
address_inb = 149;
data_ina = 16'h37f;
data_inb = 16'hf9c1;
#10;
address_ina = 150;
address_inb = 151;
data_ina = 16'hfcb6;
data_inb = 16'hfee7;
#10;
address_ina = 152;
address_inb = 153;
data_ina = 16'h347;
data_inb = 16'h158;
#10;
address_ina = 154;
address_inb = 155;
data_ina = 16'h272;
data_inb = 16'hfabf;
#10;
address_ina = 156;
address_inb = 157;
data_ina = 16'h422;
data_inb = 16'h113;
#10;
address_ina = 158;
address_inb = 159;
data_ina = 16'h5f8;
data_inb = 16'hfe3f;
#10;
address_ina = 160;
address_inb = 161;
data_ina = 16'hfd4c;
data_inb = 16'hf9cd;
#10;
address_ina = 162;
address_inb = 163;
data_ina = 16'hfcfc;
data_inb = 16'hfe9e;
#10;
address_ina = 164;
address_inb = 165;
data_ina = 16'h67c;
data_inb = 16'hfe5f;
#10;
address_ina = 166;
address_inb = 167;
data_ina = 16'h64b;
data_inb = 16'h306;
#10;
address_ina = 168;
address_inb = 169;
data_ina = 16'hfb39;
data_inb = 16'h3f7;
#10;
address_ina = 170;
address_inb = 171;
data_ina = 16'hfe38;
data_inb = 16'h89;
#10;
address_ina = 172;
address_inb = 173;
data_ina = 16'hfd1d;
data_inb = 16'hfdfe;
#10;
address_ina = 174;
address_inb = 175;
data_ina = 16'h1b8;
data_inb = 16'hfa1e;
#10;
address_ina = 176;
address_inb = 177;
data_ina = 16'hfac6;
data_inb = 16'hfc4a;
#10;
address_ina = 178;
address_inb = 179;
data_ina = 16'h61c;
data_inb = 16'hf99f;
#10;
address_ina = 180;
address_inb = 181;
data_ina = 16'h4b2;
data_inb = 16'hf9e4;
#10;
address_ina = 182;
address_inb = 183;
data_ina = 16'h2ae;
data_inb = 16'h50;
#10;
address_ina = 184;
address_inb = 185;
data_ina = 16'hff4d;
data_inb = 16'hfa5b;
#10;
address_ina = 186;
address_inb = 187;
data_ina = 16'hfde2;
data_inb = 16'hfa8a;
#10;
address_ina = 188;
address_inb = 189;
data_ina = 16'hfb5c;
data_inb = 16'h166;
#10;
address_ina = 190;
address_inb = 191;
data_ina = 16'hfe1a;
data_inb = 16'hfe57;
#10;
address_ina = 192;
address_inb = 193;
data_ina = 16'hfd4d;
data_inb = 16'hfb72;
#10;
address_ina = 194;
address_inb = 195;
data_ina = 16'hf9b0;
data_inb = 16'hfe72;
#10;
address_ina = 196;
address_inb = 197;
data_ina = 16'h547;
data_inb = 16'hfb69;
#10;
address_ina = 198;
address_inb = 199;
data_ina = 16'h475;
data_inb = 16'hfc4d;
#10;
address_ina = 200;
address_inb = 201;
data_ina = 16'hfa65;
data_inb = 16'hfc20;
#10;
address_ina = 202;
address_inb = 203;
data_ina = 16'h357;
data_inb = 16'hfdea;
#10;
address_ina = 204;
address_inb = 205;
data_ina = 16'h422;
data_inb = 16'h4cb;
#10;
address_ina = 206;
address_inb = 207;
data_ina = 16'h54f;
data_inb = 16'hfe26;
#10;
address_ina = 208;
address_inb = 209;
data_ina = 16'h170;
data_inb = 16'h18f;
#10;
address_ina = 210;
address_inb = 211;
data_ina = 16'hfe0e;
data_inb = 16'h20f;
#10;
address_ina = 212;
address_inb = 213;
data_ina = 16'h57e;
data_inb = 16'hff0f;
#10;
address_ina = 214;
address_inb = 215;
data_ina = 16'hfba2;
data_inb = 16'h338;
#10;
address_ina = 216;
address_inb = 217;
data_ina = 16'hfebc;
data_inb = 16'h2c0;
#10;
address_ina = 218;
address_inb = 219;
data_ina = 16'h5b6;
data_inb = 16'h27e;
#10;
address_ina = 220;
address_inb = 221;
data_ina = 16'h413;
data_inb = 16'h5a;
#10;
address_ina = 222;
address_inb = 223;
data_ina = 16'hfe71;
data_inb = 16'h4bf;
#10;
address_ina = 224;
address_inb = 225;
data_ina = 16'hfcc6;
data_inb = 16'hfb0d;
#10;
address_ina = 226;
address_inb = 227;
data_ina = 16'hfb0b;
data_inb = 16'h662;
#10;
address_ina = 228;
address_inb = 229;
data_ina = 16'hfb66;
data_inb = 16'h174;
#10;
address_ina = 230;
address_inb = 231;
data_ina = 16'h103;
data_inb = 16'hff12;
#10;
address_ina = 232;
address_inb = 233;
data_ina = 16'h2ac;
data_inb = 16'h77;
#10;
address_ina = 234;
address_inb = 235;
data_ina = 16'hfb92;
data_inb = 16'hfcbb;
#10;
address_ina = 236;
address_inb = 237;
data_ina = 16'h4bf;
data_inb = 16'h443;
#10;
address_ina = 238;
address_inb = 239;
data_ina = 16'hfd95;
data_inb = 16'hfb4c;
#10;
address_ina = 240;
address_inb = 241;
data_ina = 16'hfacd;
data_inb = 16'hffd6;
#10;
address_ina = 242;
address_inb = 243;
data_ina = 16'hfce0;
data_inb = 16'hfe69;
#10;
address_ina = 244;
address_inb = 245;
data_ina = 16'h2bc;
data_inb = 16'hfe32;
#10;
address_ina = 246;
address_inb = 247;
data_ina = 16'h41a;
data_inb = 16'h8d;
#10;
address_ina = 248;
address_inb = 249;
data_ina = 16'h4c5;
data_inb = 16'hfc53;
#10;
address_ina = 250;
address_inb = 251;
data_ina = 16'h108;
data_inb = 16'hfdd5;
#10;
address_ina = 252;
address_inb = 253;
data_ina = 16'hfad7;
data_inb = 16'hfece;
#10;
address_ina = 254;
address_inb = 255;
data_ina = 16'hfd93;
data_inb = 16'hff72;
#10;
        wait(init_done);
        #30
        we = 0;
        // Start processing
         
		  #38000

        start = 0;



//        wait (wr_req);
//		  wait (!wr_req);
//		   rd_req = 1;
		  wait(done);
		  #20000
rd_req = 1;
        #70 
		  start = 1;
		 #80 
wait(rd_empty)
rd_req = 0;

$display("Finished the NTT test Number %d",test_num);
////Begin test number #12//////////////
rst = 1;

//#1000
start = 1;
mode = 0; //NTT 0 // INTT 1

// Reset for a few clock cycles

#1000

rst = 0;
test_num = test_num + 1;
#1000
we = 1;
address_ina = 0;
address_inb = 1;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 2;
address_inb = 3;
data_ina = 16'h2;
data_inb = 16'hffff;
#10;
address_ina = 4;
address_inb = 5;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 6;
address_inb = 7;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 8;
address_inb = 9;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 10;
address_inb = 11;
data_ina = 16'hfffe;
data_inb = 16'h1;
#10;
address_ina = 12;
address_inb = 13;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 14;
address_inb = 15;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 16;
address_inb = 17;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 18;
address_inb = 19;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 20;
address_inb = 21;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 22;
address_inb = 23;
data_ina = 16'h0;
data_inb = 16'h2;
#10;
address_ina = 24;
address_inb = 25;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 26;
address_inb = 27;
data_ina = 16'h0;
data_inb = 16'h2;
#10;
address_ina = 28;
address_inb = 29;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 30;
address_inb = 31;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 32;
address_inb = 33;
data_ina = 16'hfffe;
data_inb = 16'hfffd;
#10;
address_ina = 34;
address_inb = 35;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 36;
address_inb = 37;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 38;
address_inb = 39;
data_ina = 16'h1;
data_inb = 16'h2;
#10;
address_ina = 40;
address_inb = 41;
data_ina = 16'h2;
data_inb = 16'h0;
#10;
address_ina = 42;
address_inb = 43;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 44;
address_inb = 45;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 46;
address_inb = 47;
data_ina = 16'h2;
data_inb = 16'hffff;
#10;
address_ina = 48;
address_inb = 49;
data_ina = 16'hfffd;
data_inb = 16'h2;
#10;
address_ina = 50;
address_inb = 51;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 52;
address_inb = 53;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 54;
address_inb = 55;
data_ina = 16'h0;
data_inb = 16'hfffe;
#10;
address_ina = 56;
address_inb = 57;
data_ina = 16'hfffe;
data_inb = 16'h0;
#10;
address_ina = 58;
address_inb = 59;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 60;
address_inb = 61;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 62;
address_inb = 63;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 64;
address_inb = 65;
data_ina = 16'hfffe;
data_inb = 16'h1;
#10;
address_ina = 66;
address_inb = 67;
data_ina = 16'hfffe;
data_inb = 16'h0;
#10;
address_ina = 68;
address_inb = 69;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 70;
address_inb = 71;
data_ina = 16'h2;
data_inb = 16'h1;
#10;
address_ina = 72;
address_inb = 73;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 74;
address_inb = 75;
data_ina = 16'h2;
data_inb = 16'h0;
#10;
address_ina = 76;
address_inb = 77;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 78;
address_inb = 79;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 80;
address_inb = 81;
data_ina = 16'hffff;
data_inb = 16'hfffe;
#10;
address_ina = 82;
address_inb = 83;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 84;
address_inb = 85;
data_ina = 16'h1;
data_inb = 16'h2;
#10;
address_ina = 86;
address_inb = 87;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 88;
address_inb = 89;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 90;
address_inb = 91;
data_ina = 16'h1;
data_inb = 16'h2;
#10;
address_ina = 92;
address_inb = 93;
data_ina = 16'h1;
data_inb = 16'hfffe;
#10;
address_ina = 94;
address_inb = 95;
data_ina = 16'h0;
data_inb = 16'hfffe;
#10;
address_ina = 96;
address_inb = 97;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 98;
address_inb = 99;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 100;
address_inb = 101;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 102;
address_inb = 103;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 104;
address_inb = 105;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 106;
address_inb = 107;
data_ina = 16'hfffe;
data_inb = 16'h2;
#10;
address_ina = 108;
address_inb = 109;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 110;
address_inb = 111;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 112;
address_inb = 113;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 114;
address_inb = 115;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 116;
address_inb = 117;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 118;
address_inb = 119;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 120;
address_inb = 121;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 122;
address_inb = 123;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 124;
address_inb = 125;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 126;
address_inb = 127;
data_ina = 16'h2;
data_inb = 16'hfffd;
#10;
address_ina = 128;
address_inb = 129;
data_ina = 16'h1;
data_inb = 16'h3;
#10;
address_ina = 130;
address_inb = 131;
data_ina = 16'h1;
data_inb = 16'h2;
#10;
address_ina = 132;
address_inb = 133;
data_ina = 16'hfffd;
data_inb = 16'h0;
#10;
address_ina = 134;
address_inb = 135;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 136;
address_inb = 137;
data_ina = 16'hfffd;
data_inb = 16'h0;
#10;
address_ina = 138;
address_inb = 139;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 140;
address_inb = 141;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 142;
address_inb = 143;
data_ina = 16'h2;
data_inb = 16'h1;
#10;
address_ina = 144;
address_inb = 145;
data_ina = 16'hfffe;
data_inb = 16'h0;
#10;
address_ina = 146;
address_inb = 147;
data_ina = 16'h1;
data_inb = 16'hfffe;
#10;
address_ina = 148;
address_inb = 149;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 150;
address_inb = 151;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 152;
address_inb = 153;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 154;
address_inb = 155;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 156;
address_inb = 157;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 158;
address_inb = 159;
data_ina = 16'h2;
data_inb = 16'hffff;
#10;
address_ina = 160;
address_inb = 161;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 162;
address_inb = 163;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 164;
address_inb = 165;
data_ina = 16'hffff;
data_inb = 16'hfffe;
#10;
address_ina = 166;
address_inb = 167;
data_ina = 16'h2;
data_inb = 16'hfffe;
#10;
address_ina = 168;
address_inb = 169;
data_ina = 16'h0;
data_inb = 16'h3;
#10;
address_ina = 170;
address_inb = 171;
data_ina = 16'h3;
data_inb = 16'hfffd;
#10;
address_ina = 172;
address_inb = 173;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 174;
address_inb = 175;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 176;
address_inb = 177;
data_ina = 16'h2;
data_inb = 16'h3;
#10;
address_ina = 178;
address_inb = 179;
data_ina = 16'h1;
data_inb = 16'h2;
#10;
address_ina = 180;
address_inb = 181;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 182;
address_inb = 183;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 184;
address_inb = 185;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 186;
address_inb = 187;
data_ina = 16'h1;
data_inb = 16'h2;
#10;
address_ina = 188;
address_inb = 189;
data_ina = 16'h2;
data_inb = 16'h1;
#10;
address_ina = 190;
address_inb = 191;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 192;
address_inb = 193;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 194;
address_inb = 195;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 196;
address_inb = 197;
data_ina = 16'h2;
data_inb = 16'hffff;
#10;
address_ina = 198;
address_inb = 199;
data_ina = 16'h0;
data_inb = 16'hfffe;
#10;
address_ina = 200;
address_inb = 201;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 202;
address_inb = 203;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 204;
address_inb = 205;
data_ina = 16'hfffe;
data_inb = 16'hfffe;
#10;
address_ina = 206;
address_inb = 207;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 208;
address_inb = 209;
data_ina = 16'hfffe;
data_inb = 16'h1;
#10;
address_ina = 210;
address_inb = 211;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 212;
address_inb = 213;
data_ina = 16'h1;
data_inb = 16'hfffe;
#10;
address_ina = 214;
address_inb = 215;
data_ina = 16'hffff;
data_inb = 16'hfffe;
#10;
address_ina = 216;
address_inb = 217;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 218;
address_inb = 219;
data_ina = 16'h0;
data_inb = 16'hfffe;
#10;
address_ina = 220;
address_inb = 221;
data_ina = 16'h2;
data_inb = 16'h3;
#10;
address_ina = 222;
address_inb = 223;
data_ina = 16'h0;
data_inb = 16'h2;
#10;
address_ina = 224;
address_inb = 225;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 226;
address_inb = 227;
data_ina = 16'hfffe;
data_inb = 16'hffff;
#10;
address_ina = 228;
address_inb = 229;
data_ina = 16'hfffd;
data_inb = 16'h0;
#10;
address_ina = 230;
address_inb = 231;
data_ina = 16'hfffe;
data_inb = 16'h2;
#10;
address_ina = 232;
address_inb = 233;
data_ina = 16'h3;
data_inb = 16'h0;
#10;
address_ina = 234;
address_inb = 235;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 236;
address_inb = 237;
data_ina = 16'hffff;
data_inb = 16'h2;
#10;
address_ina = 238;
address_inb = 239;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 240;
address_inb = 241;
data_ina = 16'h2;
data_inb = 16'h0;
#10;
address_ina = 242;
address_inb = 243;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 244;
address_inb = 245;
data_ina = 16'h2;
data_inb = 16'hffff;
#10;
address_ina = 246;
address_inb = 247;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 248;
address_inb = 249;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 250;
address_inb = 251;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 252;
address_inb = 253;
data_ina = 16'h2;
data_inb = 16'h0;
#10;
address_ina = 254;
address_inb = 255;
data_ina = 16'h0;
data_inb = 16'h3;
#10;
        wait(init_done);
        #30
        we = 0;
        // Start processing
         
		  #38000

        start = 0;



//        wait (wr_req);
//		  wait (!wr_req);
//		   rd_req = 1;
		  wait(done);
		  #20000
rd_req = 1;
        #70 
		  start = 1;
		 #80 
wait(rd_empty)
rd_req = 0;

$display("Finished the NTT test Number %d",test_num);
////Begin test number #13//////////////
rst = 1;

//#1000
start = 1;
mode = 0; //NTT 0 // INTT 1

// Reset for a few clock cycles

#1000

rst = 0;
test_num = test_num + 1;
#1000
we = 1;
address_ina = 0;
address_inb = 1;
data_ina = 16'h2;
data_inb = 16'h1;
#10;
address_ina = 2;
address_inb = 3;
data_ina = 16'hfffe;
data_inb = 16'hffff;
#10;
address_ina = 4;
address_inb = 5;
data_ina = 16'h2;
data_inb = 16'h1;
#10;
address_ina = 6;
address_inb = 7;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 8;
address_inb = 9;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 10;
address_inb = 11;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 12;
address_inb = 13;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 14;
address_inb = 15;
data_ina = 16'h1;
data_inb = 16'hfffe;
#10;
address_ina = 16;
address_inb = 17;
data_ina = 16'h2;
data_inb = 16'hfffe;
#10;
address_ina = 18;
address_inb = 19;
data_ina = 16'hfffe;
data_inb = 16'h1;
#10;
address_ina = 20;
address_inb = 21;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 22;
address_inb = 23;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 24;
address_inb = 25;
data_ina = 16'h0;
data_inb = 16'hfffe;
#10;
address_ina = 26;
address_inb = 27;
data_ina = 16'h2;
data_inb = 16'hffff;
#10;
address_ina = 28;
address_inb = 29;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 30;
address_inb = 31;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 32;
address_inb = 33;
data_ina = 16'h2;
data_inb = 16'hffff;
#10;
address_ina = 34;
address_inb = 35;
data_ina = 16'h2;
data_inb = 16'h1;
#10;
address_ina = 36;
address_inb = 37;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 38;
address_inb = 39;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 40;
address_inb = 41;
data_ina = 16'hfffe;
data_inb = 16'h0;
#10;
address_ina = 42;
address_inb = 43;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 44;
address_inb = 45;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 46;
address_inb = 47;
data_ina = 16'hfffe;
data_inb = 16'h1;
#10;
address_ina = 48;
address_inb = 49;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 50;
address_inb = 51;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 52;
address_inb = 53;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 54;
address_inb = 55;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 56;
address_inb = 57;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 58;
address_inb = 59;
data_ina = 16'h2;
data_inb = 16'h0;
#10;
address_ina = 60;
address_inb = 61;
data_ina = 16'h2;
data_inb = 16'h0;
#10;
address_ina = 62;
address_inb = 63;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 64;
address_inb = 65;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 66;
address_inb = 67;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 68;
address_inb = 69;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 70;
address_inb = 71;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 72;
address_inb = 73;
data_ina = 16'hfffe;
data_inb = 16'h1;
#10;
address_ina = 74;
address_inb = 75;
data_ina = 16'hfffd;
data_inb = 16'hffff;
#10;
address_ina = 76;
address_inb = 77;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 78;
address_inb = 79;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 80;
address_inb = 81;
data_ina = 16'h3;
data_inb = 16'h1;
#10;
address_ina = 82;
address_inb = 83;
data_ina = 16'h0;
data_inb = 16'h2;
#10;
address_ina = 84;
address_inb = 85;
data_ina = 16'h1;
data_inb = 16'h2;
#10;
address_ina = 86;
address_inb = 87;
data_ina = 16'hfffe;
data_inb = 16'h1;
#10;
address_ina = 88;
address_inb = 89;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 90;
address_inb = 91;
data_ina = 16'hfffe;
data_inb = 16'hffff;
#10;
address_ina = 92;
address_inb = 93;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 94;
address_inb = 95;
data_ina = 16'h0;
data_inb = 16'hfffe;
#10;
address_ina = 96;
address_inb = 97;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 98;
address_inb = 99;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 100;
address_inb = 101;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 102;
address_inb = 103;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 104;
address_inb = 105;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 106;
address_inb = 107;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 108;
address_inb = 109;
data_ina = 16'hfffd;
data_inb = 16'h0;
#10;
address_ina = 110;
address_inb = 111;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 112;
address_inb = 113;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 114;
address_inb = 115;
data_ina = 16'h1;
data_inb = 16'hfffe;
#10;
address_ina = 116;
address_inb = 117;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 118;
address_inb = 119;
data_ina = 16'hfffe;
data_inb = 16'hffff;
#10;
address_ina = 120;
address_inb = 121;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 122;
address_inb = 123;
data_ina = 16'hfffe;
data_inb = 16'h0;
#10;
address_ina = 124;
address_inb = 125;
data_ina = 16'h2;
data_inb = 16'h0;
#10;
address_ina = 126;
address_inb = 127;
data_ina = 16'h0;
data_inb = 16'hfffe;
#10;
address_ina = 128;
address_inb = 129;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 130;
address_inb = 131;
data_ina = 16'hfffe;
data_inb = 16'hffff;
#10;
address_ina = 132;
address_inb = 133;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 134;
address_inb = 135;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 136;
address_inb = 137;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 138;
address_inb = 139;
data_ina = 16'h1;
data_inb = 16'hfffd;
#10;
address_ina = 140;
address_inb = 141;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 142;
address_inb = 143;
data_ina = 16'h2;
data_inb = 16'h1;
#10;
address_ina = 144;
address_inb = 145;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 146;
address_inb = 147;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 148;
address_inb = 149;
data_ina = 16'h0;
data_inb = 16'hfffe;
#10;
address_ina = 150;
address_inb = 151;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 152;
address_inb = 153;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 154;
address_inb = 155;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 156;
address_inb = 157;
data_ina = 16'h0;
data_inb = 16'hfffe;
#10;
address_ina = 158;
address_inb = 159;
data_ina = 16'hffff;
data_inb = 16'hfffe;
#10;
address_ina = 160;
address_inb = 161;
data_ina = 16'h0;
data_inb = 16'h2;
#10;
address_ina = 162;
address_inb = 163;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 164;
address_inb = 165;
data_ina = 16'h2;
data_inb = 16'hfffd;
#10;
address_ina = 166;
address_inb = 167;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 168;
address_inb = 169;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 170;
address_inb = 171;
data_ina = 16'hfffe;
data_inb = 16'h1;
#10;
address_ina = 172;
address_inb = 173;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 174;
address_inb = 175;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 176;
address_inb = 177;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 178;
address_inb = 179;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 180;
address_inb = 181;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 182;
address_inb = 183;
data_ina = 16'hffff;
data_inb = 16'hfffe;
#10;
address_ina = 184;
address_inb = 185;
data_ina = 16'h0;
data_inb = 16'hfffe;
#10;
address_ina = 186;
address_inb = 187;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 188;
address_inb = 189;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 190;
address_inb = 191;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 192;
address_inb = 193;
data_ina = 16'h2;
data_inb = 16'h1;
#10;
address_ina = 194;
address_inb = 195;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 196;
address_inb = 197;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 198;
address_inb = 199;
data_ina = 16'hfffe;
data_inb = 16'h1;
#10;
address_ina = 200;
address_inb = 201;
data_ina = 16'hffff;
data_inb = 16'hfffe;
#10;
address_ina = 202;
address_inb = 203;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 204;
address_inb = 205;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 206;
address_inb = 207;
data_ina = 16'hfffe;
data_inb = 16'hffff;
#10;
address_ina = 208;
address_inb = 209;
data_ina = 16'hfffe;
data_inb = 16'h0;
#10;
address_ina = 210;
address_inb = 211;
data_ina = 16'hfffe;
data_inb = 16'hfffe;
#10;
address_ina = 212;
address_inb = 213;
data_ina = 16'hfffe;
data_inb = 16'h1;
#10;
address_ina = 214;
address_inb = 215;
data_ina = 16'h2;
data_inb = 16'h1;
#10;
address_ina = 216;
address_inb = 217;
data_ina = 16'h2;
data_inb = 16'hffff;
#10;
address_ina = 218;
address_inb = 219;
data_ina = 16'hffff;
data_inb = 16'hfffe;
#10;
address_ina = 220;
address_inb = 221;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 222;
address_inb = 223;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 224;
address_inb = 225;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 226;
address_inb = 227;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 228;
address_inb = 229;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 230;
address_inb = 231;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 232;
address_inb = 233;
data_ina = 16'h0;
data_inb = 16'h2;
#10;
address_ina = 234;
address_inb = 235;
data_ina = 16'h0;
data_inb = 16'h3;
#10;
address_ina = 236;
address_inb = 237;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 238;
address_inb = 239;
data_ina = 16'h1;
data_inb = 16'hfffe;
#10;
address_ina = 240;
address_inb = 241;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 242;
address_inb = 243;
data_ina = 16'hfffe;
data_inb = 16'hffff;
#10;
address_ina = 244;
address_inb = 245;
data_ina = 16'h0;
data_inb = 16'h2;
#10;
address_ina = 246;
address_inb = 247;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 248;
address_inb = 249;
data_ina = 16'hffff;
data_inb = 16'h3;
#10;
address_ina = 250;
address_inb = 251;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 252;
address_inb = 253;
data_ina = 16'h0;
data_inb = 16'hfffe;
#10;
address_ina = 254;
address_inb = 255;
data_ina = 16'h3;
data_inb = 16'h1;
#10;
        wait(init_done);
        #30
        we = 0;
        // Start processing
         
		  #38000

        start = 0;



//        wait (wr_req);
//		  wait (!wr_req);
//		   rd_req = 1;
		  wait(done);
		  #20000
rd_req = 1;
        #70 
		  start = 1;
		 #80 
wait(rd_empty)
rd_req = 0;

$display("Finished the NTT test Number %d",test_num);
////Begin test number #14//////////////
rst = 1;

//#1000
start = 1;
mode = 1; //NTT 0 // INTT 1

// Reset for a few clock cycles

#1000

rst = 0;
test_num = test_num + 1;
#1000
we = 1;
address_ina = 0;
address_inb = 1;
data_ina = 16'h410;
data_inb = 16'hf9e2;
#10;
address_ina = 2;
address_inb = 3;
data_ina = 16'h3be;
data_inb = 16'h43e;
#10;
address_ina = 4;
address_inb = 5;
data_ina = 16'h321;
data_inb = 16'h3f2;
#10;
address_ina = 6;
address_inb = 7;
data_ina = 16'hfac5;
data_inb = 16'h255;
#10;
address_ina = 8;
address_inb = 9;
data_ina = 16'hfe2b;
data_inb = 16'hff3d;
#10;
address_ina = 10;
address_inb = 11;
data_ina = 16'h420;
data_inb = 16'hfec1;
#10;
address_ina = 12;
address_inb = 13;
data_ina = 16'h215;
data_inb = 16'hfebe;
#10;
address_ina = 14;
address_inb = 15;
data_ina = 16'hfa07;
data_inb = 16'hfb98;
#10;
address_ina = 16;
address_inb = 17;
data_ina = 16'hff9a;
data_inb = 16'h41c;
#10;
address_ina = 18;
address_inb = 19;
data_ina = 16'hfcc0;
data_inb = 16'h17;
#10;
address_ina = 20;
address_inb = 21;
data_ina = 16'hfab0;
data_inb = 16'h2d8;
#10;
address_ina = 22;
address_inb = 23;
data_ina = 16'h2e3;
data_inb = 16'h665;
#10;
address_ina = 24;
address_inb = 25;
data_ina = 16'hfd2b;
data_inb = 16'h394;
#10;
address_ina = 26;
address_inb = 27;
data_ina = 16'hf98e;
data_inb = 16'h23c;
#10;
address_ina = 28;
address_inb = 29;
data_ina = 16'h560;
data_inb = 16'h313;
#10;
address_ina = 30;
address_inb = 31;
data_ina = 16'h203;
data_inb = 16'hfcd1;
#10;
address_ina = 32;
address_inb = 33;
data_ina = 16'h634;
data_inb = 16'hffcc;
#10;
address_ina = 34;
address_inb = 35;
data_ina = 16'hfeb6;
data_inb = 16'hfcc7;
#10;
address_ina = 36;
address_inb = 37;
data_ina = 16'hfa06;
data_inb = 16'hf98d;
#10;
address_ina = 38;
address_inb = 39;
data_ina = 16'h5fe;
data_inb = 16'hfcc4;
#10;
address_ina = 40;
address_inb = 41;
data_ina = 16'hfec6;
data_inb = 16'hfadd;
#10;
address_ina = 42;
address_inb = 43;
data_ina = 16'h92;
data_inb = 16'h25e;
#10;
address_ina = 44;
address_inb = 45;
data_ina = 16'h203;
data_inb = 16'hfbea;
#10;
address_ina = 46;
address_inb = 47;
data_ina = 16'h1b7;
data_inb = 16'hfc35;
#10;
address_ina = 48;
address_inb = 49;
data_ina = 16'h2db;
data_inb = 16'h156;
#10;
address_ina = 50;
address_inb = 51;
data_ina = 16'h4d5;
data_inb = 16'h40;
#10;
address_ina = 52;
address_inb = 53;
data_ina = 16'h1b;
data_inb = 16'hff7a;
#10;
address_ina = 54;
address_inb = 55;
data_ina = 16'h366;
data_inb = 16'hfa55;
#10;
address_ina = 56;
address_inb = 57;
data_ina = 16'h29c;
data_inb = 16'hfd96;
#10;
address_ina = 58;
address_inb = 59;
data_ina = 16'h515;
data_inb = 16'hfcd3;
#10;
address_ina = 60;
address_inb = 61;
data_ina = 16'h341;
data_inb = 16'h3ed;
#10;
address_ina = 62;
address_inb = 63;
data_ina = 16'h2e5;
data_inb = 16'h5a2;
#10;
address_ina = 64;
address_inb = 65;
data_ina = 16'h1e0;
data_inb = 16'hf9e3;
#10;
address_ina = 66;
address_inb = 67;
data_ina = 16'hfd01;
data_inb = 16'h262;
#10;
address_ina = 68;
address_inb = 69;
data_ina = 16'h42d;
data_inb = 16'hffed;
#10;
address_ina = 70;
address_inb = 71;
data_ina = 16'hfa45;
data_inb = 16'h2dd;
#10;
address_ina = 72;
address_inb = 73;
data_ina = 16'hffac;
data_inb = 16'h2a;
#10;
address_ina = 74;
address_inb = 75;
data_ina = 16'hfd4d;
data_inb = 16'h5a8;
#10;
address_ina = 76;
address_inb = 77;
data_ina = 16'hfd9c;
data_inb = 16'hff36;
#10;
address_ina = 78;
address_inb = 79;
data_ina = 16'h158;
data_inb = 16'hfbf3;
#10;
address_ina = 80;
address_inb = 81;
data_ina = 16'h676;
data_inb = 16'hfb11;
#10;
address_ina = 82;
address_inb = 83;
data_ina = 16'hfbd0;
data_inb = 16'h235;
#10;
address_ina = 84;
address_inb = 85;
data_ina = 16'h354;
data_inb = 16'h74;
#10;
address_ina = 86;
address_inb = 87;
data_ina = 16'hfdf7;
data_inb = 16'hfa56;
#10;
address_ina = 88;
address_inb = 89;
data_ina = 16'hfc60;
data_inb = 16'hfa5d;
#10;
address_ina = 90;
address_inb = 91;
data_ina = 16'hfddd;
data_inb = 16'h37f;
#10;
address_ina = 92;
address_inb = 93;
data_ina = 16'hff80;
data_inb = 16'hfba5;
#10;
address_ina = 94;
address_inb = 95;
data_ina = 16'h4c3;
data_inb = 16'hfa4c;
#10;
address_ina = 96;
address_inb = 97;
data_ina = 16'h51b;
data_inb = 16'hfe6d;
#10;
address_ina = 98;
address_inb = 99;
data_ina = 16'h53f;
data_inb = 16'hfe1c;
#10;
address_ina = 100;
address_inb = 101;
data_ina = 16'h1a0;
data_inb = 16'hf9fb;
#10;
address_ina = 102;
address_inb = 103;
data_ina = 16'h5b;
data_inb = 16'hfdb7;
#10;
address_ina = 104;
address_inb = 105;
data_ina = 16'ha3;
data_inb = 16'h3bc;
#10;
address_ina = 106;
address_inb = 107;
data_ina = 16'hfe2b;
data_inb = 16'hf9a5;
#10;
address_ina = 108;
address_inb = 109;
data_ina = 16'hfa79;
data_inb = 16'h4cd;
#10;
address_ina = 110;
address_inb = 111;
data_ina = 16'hfaac;
data_inb = 16'hfce2;
#10;
address_ina = 112;
address_inb = 113;
data_ina = 16'hfabb;
data_inb = 16'hfa83;
#10;
address_ina = 114;
address_inb = 115;
data_ina = 16'h124;
data_inb = 16'hfb1b;
#10;
address_ina = 116;
address_inb = 117;
data_ina = 16'hfe3d;
data_inb = 16'h65d;
#10;
address_ina = 118;
address_inb = 119;
data_ina = 16'h15d;
data_inb = 16'hff55;
#10;
address_ina = 120;
address_inb = 121;
data_ina = 16'h1ac;
data_inb = 16'hf4;
#10;
address_ina = 122;
address_inb = 123;
data_ina = 16'hfac2;
data_inb = 16'hee;
#10;
address_ina = 124;
address_inb = 125;
data_ina = 16'hfd7c;
data_inb = 16'h528;
#10;
address_ina = 126;
address_inb = 127;
data_ina = 16'hbc;
data_inb = 16'h17c;
#10;
address_ina = 128;
address_inb = 129;
data_ina = 16'h5e6;
data_inb = 16'hfb05;
#10;
address_ina = 130;
address_inb = 131;
data_ina = 16'h481;
data_inb = 16'h232;
#10;
address_ina = 132;
address_inb = 133;
data_ina = 16'hfc80;
data_inb = 16'hfdd3;
#10;
address_ina = 134;
address_inb = 135;
data_ina = 16'h6a;
data_inb = 16'h21f;
#10;
address_ina = 136;
address_inb = 137;
data_ina = 16'h5e5;
data_inb = 16'h1ff;
#10;
address_ina = 138;
address_inb = 139;
data_ina = 16'h377;
data_inb = 16'hfc81;
#10;
address_ina = 140;
address_inb = 141;
data_ina = 16'hfabe;
data_inb = 16'hfd73;
#10;
address_ina = 142;
address_inb = 143;
data_ina = 16'h5e;
data_inb = 16'he7;
#10;
address_ina = 144;
address_inb = 145;
data_ina = 16'h562;
data_inb = 16'h8;
#10;
address_ina = 146;
address_inb = 147;
data_ina = 16'h40a;
data_inb = 16'h9c;
#10;
address_ina = 148;
address_inb = 149;
data_ina = 16'h7;
data_inb = 16'h5ef;
#10;
address_ina = 150;
address_inb = 151;
data_ina = 16'hfbdd;
data_inb = 16'hfb00;
#10;
address_ina = 152;
address_inb = 153;
data_ina = 16'hfd29;
data_inb = 16'hfa94;
#10;
address_ina = 154;
address_inb = 155;
data_ina = 16'h134;
data_inb = 16'hfe63;
#10;
address_ina = 156;
address_inb = 157;
data_ina = 16'hfeb0;
data_inb = 16'h401;
#10;
address_ina = 158;
address_inb = 159;
data_ina = 16'hfb33;
data_inb = 16'hf9be;
#10;
address_ina = 160;
address_inb = 161;
data_ina = 16'h2fc;
data_inb = 16'hffdd;
#10;
address_ina = 162;
address_inb = 163;
data_ina = 16'hfb4d;
data_inb = 16'hfaf5;
#10;
address_ina = 164;
address_inb = 165;
data_ina = 16'h11e;
data_inb = 16'h1c5;
#10;
address_ina = 166;
address_inb = 167;
data_ina = 16'hfae6;
data_inb = 16'hc6;
#10;
address_ina = 168;
address_inb = 169;
data_ina = 16'hfd4e;
data_inb = 16'hfae6;
#10;
address_ina = 170;
address_inb = 171;
data_ina = 16'h35f;
data_inb = 16'h25b;
#10;
address_ina = 172;
address_inb = 173;
data_ina = 16'h2db;
data_inb = 16'h10c;
#10;
address_ina = 174;
address_inb = 175;
data_ina = 16'hfb6c;
data_inb = 16'hfa91;
#10;
address_ina = 176;
address_inb = 177;
data_ina = 16'h17d;
data_inb = 16'hfbbd;
#10;
address_ina = 178;
address_inb = 179;
data_ina = 16'h8c;
data_inb = 16'hff60;
#10;
address_ina = 180;
address_inb = 181;
data_ina = 16'hf9ea;
data_inb = 16'h620;
#10;
address_ina = 182;
address_inb = 183;
data_ina = 16'h1d1;
data_inb = 16'h22c;
#10;
address_ina = 184;
address_inb = 185;
data_ina = 16'h2a7;
data_inb = 16'h66;
#10;
address_ina = 186;
address_inb = 187;
data_ina = 16'hffd2;
data_inb = 16'hfc6b;
#10;
address_ina = 188;
address_inb = 189;
data_ina = 16'hff84;
data_inb = 16'hfcec;
#10;
address_ina = 190;
address_inb = 191;
data_ina = 16'h447;
data_inb = 16'hfa93;
#10;
address_ina = 192;
address_inb = 193;
data_ina = 16'h412;
data_inb = 16'hfae7;
#10;
address_ina = 194;
address_inb = 195;
data_ina = 16'hfb10;
data_inb = 16'hfc21;
#10;
address_ina = 196;
address_inb = 197;
data_ina = 16'h323;
data_inb = 16'h649;
#10;
address_ina = 198;
address_inb = 199;
data_ina = 16'hfee4;
data_inb = 16'hfeb5;
#10;
address_ina = 200;
address_inb = 201;
data_ina = 16'h441;
data_inb = 16'h21a;
#10;
address_ina = 202;
address_inb = 203;
data_ina = 16'h395;
data_inb = 16'heb;
#10;
address_ina = 204;
address_inb = 205;
data_ina = 16'hfca3;
data_inb = 16'h2f0;
#10;
address_ina = 206;
address_inb = 207;
data_ina = 16'h593;
data_inb = 16'hfa36;
#10;
address_ina = 208;
address_inb = 209;
data_ina = 16'hfac5;
data_inb = 16'hff18;
#10;
address_ina = 210;
address_inb = 211;
data_ina = 16'h288;
data_inb = 16'hfe04;
#10;
address_ina = 212;
address_inb = 213;
data_ina = 16'hfb92;
data_inb = 16'hfe33;
#10;
address_ina = 214;
address_inb = 215;
data_ina = 16'hfaad;
data_inb = 16'hfb26;
#10;
address_ina = 216;
address_inb = 217;
data_ina = 16'hff11;
data_inb = 16'hfb40;
#10;
address_ina = 218;
address_inb = 219;
data_ina = 16'h38;
data_inb = 16'hfa68;
#10;
address_ina = 220;
address_inb = 221;
data_ina = 16'hfd12;
data_inb = 16'hfa27;
#10;
address_ina = 222;
address_inb = 223;
data_ina = 16'h4e1;
data_inb = 16'h3e5;
#10;
address_ina = 224;
address_inb = 225;
data_ina = 16'hf990;
data_inb = 16'h317;
#10;
address_ina = 226;
address_inb = 227;
data_ina = 16'hf98e;
data_inb = 16'h53f;
#10;
address_ina = 228;
address_inb = 229;
data_ina = 16'hfa55;
data_inb = 16'h524;
#10;
address_ina = 230;
address_inb = 231;
data_ina = 16'hfd77;
data_inb = 16'h7;
#10;
address_ina = 232;
address_inb = 233;
data_ina = 16'hfe84;
data_inb = 16'h212;
#10;
address_ina = 234;
address_inb = 235;
data_ina = 16'hfbe2;
data_inb = 16'hfd33;
#10;
address_ina = 236;
address_inb = 237;
data_ina = 16'hfde4;
data_inb = 16'h98;
#10;
address_ina = 238;
address_inb = 239;
data_ina = 16'hfc36;
data_inb = 16'hfd85;
#10;
address_ina = 240;
address_inb = 241;
data_ina = 16'h325;
data_inb = 16'h37a;
#10;
address_ina = 242;
address_inb = 243;
data_ina = 16'hfa98;
data_inb = 16'hfbcb;
#10;
address_ina = 244;
address_inb = 245;
data_ina = 16'h12c;
data_inb = 16'h33f;
#10;
address_ina = 246;
address_inb = 247;
data_ina = 16'hfcde;
data_inb = 16'h407;
#10;
address_ina = 248;
address_inb = 249;
data_ina = 16'h520;
data_inb = 16'hfb70;
#10;
address_ina = 250;
address_inb = 251;
data_ina = 16'hff95;
data_inb = 16'h5e6;
#10;
address_ina = 252;
address_inb = 253;
data_ina = 16'hff84;
data_inb = 16'h166;
#10;
address_ina = 254;
address_inb = 255;
data_ina = 16'h66b;
data_inb = 16'h477;
#10;
        wait(init_done);
        #30
        we = 0;
        // Start processing
         
		  #38000

        start = 0;



//        wait (wr_req);
//		  wait (!wr_req);
//		   rd_req = 1;
		  wait(done);
		  #20000
rd_req = 1;
        #70 
		  start = 1;
		 #80 
wait(rd_empty)
rd_req = 0;

$display("Finished the NTT test Number %d",test_num);
////Begin test number #15//////////////
rst = 1;

//#1000
start = 1;
mode = 1; //NTT 0 // INTT 1

// Reset for a few clock cycles

#1000

rst = 0;
test_num = test_num + 1;
#1000
we = 1;
address_ina = 0;
address_inb = 1;
data_ina = 16'hfe35;
data_inb = 16'h378;
#10;
address_ina = 2;
address_inb = 3;
data_ina = 16'h455;
data_inb = 16'hfed6;
#10;
address_ina = 4;
address_inb = 5;
data_ina = 16'h62e;
data_inb = 16'hfaec;
#10;
address_ina = 6;
address_inb = 7;
data_ina = 16'hfe8d;
data_inb = 16'hfe7f;
#10;
address_ina = 8;
address_inb = 9;
data_ina = 16'hfe97;
data_inb = 16'hfbac;
#10;
address_ina = 10;
address_inb = 11;
data_ina = 16'hf9eb;
data_inb = 16'h65a;
#10;
address_ina = 12;
address_inb = 13;
data_ina = 16'hfd5b;
data_inb = 16'h57;
#10;
address_ina = 14;
address_inb = 15;
data_ina = 16'h460;
data_inb = 16'hf9ae;
#10;
address_ina = 16;
address_inb = 17;
data_ina = 16'h217;
data_inb = 16'h28a;
#10;
address_ina = 18;
address_inb = 19;
data_ina = 16'h436;
data_inb = 16'h36d;
#10;
address_ina = 20;
address_inb = 21;
data_ina = 16'h594;
data_inb = 16'h5d6;
#10;
address_ina = 22;
address_inb = 23;
data_ina = 16'hff50;
data_inb = 16'h1e0;
#10;
address_ina = 24;
address_inb = 25;
data_ina = 16'hfe0a;
data_inb = 16'hfdc3;
#10;
address_ina = 26;
address_inb = 27;
data_ina = 16'hfe7a;
data_inb = 16'hf9f3;
#10;
address_ina = 28;
address_inb = 29;
data_ina = 16'hfa10;
data_inb = 16'hf9b3;
#10;
address_ina = 30;
address_inb = 31;
data_ina = 16'hfa4a;
data_inb = 16'h2b8;
#10;
address_ina = 32;
address_inb = 33;
data_ina = 16'hff93;
data_inb = 16'hfe15;
#10;
address_ina = 34;
address_inb = 35;
data_ina = 16'h271;
data_inb = 16'hf9bf;
#10;
address_ina = 36;
address_inb = 37;
data_ina = 16'h579;
data_inb = 16'hff02;
#10;
address_ina = 38;
address_inb = 39;
data_ina = 16'h47e;
data_inb = 16'hfaed;
#10;
address_ina = 40;
address_inb = 41;
data_ina = 16'h548;
data_inb = 16'h427;
#10;
address_ina = 42;
address_inb = 43;
data_ina = 16'h1ac;
data_inb = 16'h608;
#10;
address_ina = 44;
address_inb = 45;
data_ina = 16'h6b;
data_inb = 16'hfcdb;
#10;
address_ina = 46;
address_inb = 47;
data_ina = 16'h1e6;
data_inb = 16'hfd4e;
#10;
address_ina = 48;
address_inb = 49;
data_ina = 16'hfe36;
data_inb = 16'hbd;
#10;
address_ina = 50;
address_inb = 51;
data_ina = 16'h42e;
data_inb = 16'h36f;
#10;
address_ina = 52;
address_inb = 53;
data_ina = 16'h3ca;
data_inb = 16'h1;
#10;
address_ina = 54;
address_inb = 55;
data_ina = 16'h473;
data_inb = 16'h5ce;
#10;
address_ina = 56;
address_inb = 57;
data_ina = 16'h79;
data_inb = 16'hf9e7;
#10;
address_ina = 58;
address_inb = 59;
data_ina = 16'hfb1d;
data_inb = 16'hff51;
#10;
address_ina = 60;
address_inb = 61;
data_ina = 16'h32c;
data_inb = 16'h4fc;
#10;
address_ina = 62;
address_inb = 63;
data_ina = 16'h8f;
data_inb = 16'hfe55;
#10;
address_ina = 64;
address_inb = 65;
data_ina = 16'h13f;
data_inb = 16'hfbe0;
#10;
address_ina = 66;
address_inb = 67;
data_ina = 16'hfc37;
data_inb = 16'h223;
#10;
address_ina = 68;
address_inb = 69;
data_ina = 16'h149;
data_inb = 16'hf2;
#10;
address_ina = 70;
address_inb = 71;
data_ina = 16'hfef9;
data_inb = 16'h2d9;
#10;
address_ina = 72;
address_inb = 73;
data_ina = 16'hfa7f;
data_inb = 16'hfc55;
#10;
address_ina = 74;
address_inb = 75;
data_ina = 16'h2c;
data_inb = 16'hfbdd;
#10;
address_ina = 76;
address_inb = 77;
data_ina = 16'hffcf;
data_inb = 16'h2b2;
#10;
address_ina = 78;
address_inb = 79;
data_ina = 16'hfdd1;
data_inb = 16'h36;
#10;
address_ina = 80;
address_inb = 81;
data_ina = 16'h27d;
data_inb = 16'hfffe;
#10;
address_ina = 82;
address_inb = 83;
data_ina = 16'h5f5;
data_inb = 16'h43b;
#10;
address_ina = 84;
address_inb = 85;
data_ina = 16'hf994;
data_inb = 16'hfa55;
#10;
address_ina = 86;
address_inb = 87;
data_ina = 16'hfd6b;
data_inb = 16'hfe50;
#10;
address_ina = 88;
address_inb = 89;
data_ina = 16'h58d;
data_inb = 16'h44f;
#10;
address_ina = 90;
address_inb = 91;
data_ina = 16'h1ad;
data_inb = 16'hfd8f;
#10;
address_ina = 92;
address_inb = 93;
data_ina = 16'hffab;
data_inb = 16'hfa0e;
#10;
address_ina = 94;
address_inb = 95;
data_ina = 16'hff5b;
data_inb = 16'h17c;
#10;
address_ina = 96;
address_inb = 97;
data_ina = 16'hfb0b;
data_inb = 16'h622;
#10;
address_ina = 98;
address_inb = 99;
data_ina = 16'hfcdc;
data_inb = 16'h1df;
#10;
address_ina = 100;
address_inb = 101;
data_ina = 16'h2e5;
data_inb = 16'hf9be;
#10;
address_ina = 102;
address_inb = 103;
data_ina = 16'h3f;
data_inb = 16'hfbb2;
#10;
address_ina = 104;
address_inb = 105;
data_ina = 16'h3ef;
data_inb = 16'h1a4;
#10;
address_ina = 106;
address_inb = 107;
data_ina = 16'hfdb6;
data_inb = 16'h4e2;
#10;
address_ina = 108;
address_inb = 109;
data_ina = 16'hfbc3;
data_inb = 16'hfbc4;
#10;
address_ina = 110;
address_inb = 111;
data_ina = 16'hfef6;
data_inb = 16'hf9ee;
#10;
address_ina = 112;
address_inb = 113;
data_ina = 16'hf9d9;
data_inb = 16'hff25;
#10;
address_ina = 114;
address_inb = 115;
data_ina = 16'hf9c1;
data_inb = 16'h275;
#10;
address_ina = 116;
address_inb = 117;
data_ina = 16'h65f;
data_inb = 16'hfa25;
#10;
address_ina = 118;
address_inb = 119;
data_ina = 16'h549;
data_inb = 16'h124;
#10;
address_ina = 120;
address_inb = 121;
data_ina = 16'h285;
data_inb = 16'h430;
#10;
address_ina = 122;
address_inb = 123;
data_ina = 16'hfebd;
data_inb = 16'hfb24;
#10;
address_ina = 124;
address_inb = 125;
data_ina = 16'hfa3a;
data_inb = 16'hfb03;
#10;
address_ina = 126;
address_inb = 127;
data_ina = 16'hfef2;
data_inb = 16'hff2c;
#10;
address_ina = 128;
address_inb = 129;
data_ina = 16'h175;
data_inb = 16'hfc8d;
#10;
address_ina = 130;
address_inb = 131;
data_ina = 16'hf7;
data_inb = 16'hfc0c;
#10;
address_ina = 132;
address_inb = 133;
data_ina = 16'hfdfb;
data_inb = 16'h49a;
#10;
address_ina = 134;
address_inb = 135;
data_ina = 16'hfffb;
data_inb = 16'h5ac;
#10;
address_ina = 136;
address_inb = 137;
data_ina = 16'hfe8a;
data_inb = 16'hff37;
#10;
address_ina = 138;
address_inb = 139;
data_ina = 16'hfd7b;
data_inb = 16'hfe98;
#10;
address_ina = 140;
address_inb = 141;
data_ina = 16'h451;
data_inb = 16'h19a;
#10;
address_ina = 142;
address_inb = 143;
data_ina = 16'h5ae;
data_inb = 16'hfdef;
#10;
address_ina = 144;
address_inb = 145;
data_ina = 16'h495;
data_inb = 16'h55;
#10;
address_ina = 146;
address_inb = 147;
data_ina = 16'hfc74;
data_inb = 16'hfb6a;
#10;
address_ina = 148;
address_inb = 149;
data_ina = 16'hfa0d;
data_inb = 16'h40d;
#10;
address_ina = 150;
address_inb = 151;
data_ina = 16'hffe6;
data_inb = 16'h51e;
#10;
address_ina = 152;
address_inb = 153;
data_ina = 16'hfd17;
data_inb = 16'hff28;
#10;
address_ina = 154;
address_inb = 155;
data_ina = 16'hfd08;
data_inb = 16'hfac1;
#10;
address_ina = 156;
address_inb = 157;
data_ina = 16'hfb44;
data_inb = 16'hfe08;
#10;
address_ina = 158;
address_inb = 159;
data_ina = 16'h57;
data_inb = 16'hfae6;
#10;
address_ina = 160;
address_inb = 161;
data_ina = 16'hfb04;
data_inb = 16'hfdb8;
#10;
address_ina = 162;
address_inb = 163;
data_ina = 16'hfe58;
data_inb = 16'h2ba;
#10;
address_ina = 164;
address_inb = 165;
data_ina = 16'hfb75;
data_inb = 16'h4ed;
#10;
address_ina = 166;
address_inb = 167;
data_ina = 16'hff1c;
data_inb = 16'hfbba;
#10;
address_ina = 168;
address_inb = 169;
data_ina = 16'h55c;
data_inb = 16'h5cf;
#10;
address_ina = 170;
address_inb = 171;
data_ina = 16'hfd7d;
data_inb = 16'hfa08;
#10;
address_ina = 172;
address_inb = 173;
data_ina = 16'hfc5e;
data_inb = 16'h4c8;
#10;
address_ina = 174;
address_inb = 175;
data_ina = 16'h6a;
data_inb = 16'h2c;
#10;
address_ina = 176;
address_inb = 177;
data_ina = 16'hfc15;
data_inb = 16'h82;
#10;
address_ina = 178;
address_inb = 179;
data_ina = 16'hfaf8;
data_inb = 16'h3ef;
#10;
address_ina = 180;
address_inb = 181;
data_ina = 16'h30e;
data_inb = 16'h507;
#10;
address_ina = 182;
address_inb = 183;
data_ina = 16'h445;
data_inb = 16'hfc77;
#10;
address_ina = 184;
address_inb = 185;
data_ina = 16'hfdd5;
data_inb = 16'h353;
#10;
address_ina = 186;
address_inb = 187;
data_ina = 16'h53d;
data_inb = 16'hfdf4;
#10;
address_ina = 188;
address_inb = 189;
data_ina = 16'hfd55;
data_inb = 16'hfa3a;
#10;
address_ina = 190;
address_inb = 191;
data_ina = 16'h1b7;
data_inb = 16'hfcaf;
#10;
address_ina = 192;
address_inb = 193;
data_ina = 16'hfb55;
data_inb = 16'hfa4b;
#10;
address_ina = 194;
address_inb = 195;
data_ina = 16'hfbe6;
data_inb = 16'hfb12;
#10;
address_ina = 196;
address_inb = 197;
data_ina = 16'h82;
data_inb = 16'h654;
#10;
address_ina = 198;
address_inb = 199;
data_ina = 16'hff49;
data_inb = 16'hff48;
#10;
address_ina = 200;
address_inb = 201;
data_ina = 16'h158;
data_inb = 16'hfb15;
#10;
address_ina = 202;
address_inb = 203;
data_ina = 16'hfa01;
data_inb = 16'h2f4;
#10;
address_ina = 204;
address_inb = 205;
data_ina = 16'h4a5;
data_inb = 16'h3f0;
#10;
address_ina = 206;
address_inb = 207;
data_ina = 16'hfd82;
data_inb = 16'h582;
#10;
address_ina = 208;
address_inb = 209;
data_ina = 16'h28f;
data_inb = 16'h4be;
#10;
address_ina = 210;
address_inb = 211;
data_ina = 16'h223;
data_inb = 16'h5be;
#10;
address_ina = 212;
address_inb = 213;
data_ina = 16'h518;
data_inb = 16'h214;
#10;
address_ina = 214;
address_inb = 215;
data_ina = 16'hfa8e;
data_inb = 16'hfca1;
#10;
address_ina = 216;
address_inb = 217;
data_ina = 16'hfafd;
data_inb = 16'hff0b;
#10;
address_ina = 218;
address_inb = 219;
data_ina = 16'h2ec;
data_inb = 16'h443;
#10;
address_ina = 220;
address_inb = 221;
data_ina = 16'h264;
data_inb = 16'h504;
#10;
address_ina = 222;
address_inb = 223;
data_ina = 16'hfb77;
data_inb = 16'hfc75;
#10;
address_ina = 224;
address_inb = 225;
data_ina = 16'hfd1a;
data_inb = 16'hfff4;
#10;
address_ina = 226;
address_inb = 227;
data_ina = 16'hfc57;
data_inb = 16'hff63;
#10;
address_ina = 228;
address_inb = 229;
data_ina = 16'h422;
data_inb = 16'h61a;
#10;
address_ina = 230;
address_inb = 231;
data_ina = 16'hfb3d;
data_inb = 16'h2e8;
#10;
address_ina = 232;
address_inb = 233;
data_ina = 16'h5a3;
data_inb = 16'hfb7a;
#10;
address_ina = 234;
address_inb = 235;
data_ina = 16'hfae8;
data_inb = 16'h57;
#10;
address_ina = 236;
address_inb = 237;
data_ina = 16'hfde6;
data_inb = 16'hf9b4;
#10;
address_ina = 238;
address_inb = 239;
data_ina = 16'h15d;
data_inb = 16'h2d2;
#10;
address_ina = 240;
address_inb = 241;
data_ina = 16'h493;
data_inb = 16'h163;
#10;
address_ina = 242;
address_inb = 243;
data_ina = 16'h322;
data_inb = 16'hffe4;
#10;
address_ina = 244;
address_inb = 245;
data_ina = 16'h466;
data_inb = 16'h144;
#10;
address_ina = 246;
address_inb = 247;
data_ina = 16'h366;
data_inb = 16'h623;
#10;
address_ina = 248;
address_inb = 249;
data_ina = 16'h48b;
data_inb = 16'h482;
#10;
address_ina = 250;
address_inb = 251;
data_ina = 16'hfb56;
data_inb = 16'h4;
#10;
address_ina = 252;
address_inb = 253;
data_ina = 16'hfeef;
data_inb = 16'h216;
#10;
address_ina = 254;
address_inb = 255;
data_ina = 16'h168;
data_inb = 16'heb;
#10;
        wait(init_done);
        #30
        we = 0;
        // Start processing
         
		  #38000

        start = 0;



//        wait (wr_req);
//		  wait (!wr_req);
//		   rd_req = 1;
		  wait(done);
		  #20000
rd_req = 1;
        #70 
		  start = 1;
		 #80 
wait(rd_empty)
rd_req = 0;

$display("Finished the NTT test Number %d",test_num);
////Begin test number #16//////////////
rst = 1;

//#1000
start = 1;
mode = 1; //NTT 0 // INTT 1

// Reset for a few clock cycles

#1000

rst = 0;
test_num = test_num + 1;
#1000
we = 1;
address_ina = 0;
address_inb = 1;
data_ina = 16'hfd21;
data_inb = 16'h277;
#10;
address_ina = 2;
address_inb = 3;
data_ina = 16'h2e1;
data_inb = 16'hfb1f;
#10;
address_ina = 4;
address_inb = 5;
data_ina = 16'h5c6;
data_inb = 16'h132;
#10;
address_ina = 6;
address_inb = 7;
data_ina = 16'h4e2;
data_inb = 16'hc1;
#10;
address_ina = 8;
address_inb = 9;
data_ina = 16'hf9cb;
data_inb = 16'hfaf0;
#10;
address_ina = 10;
address_inb = 11;
data_ina = 16'hfef0;
data_inb = 16'hff0c;
#10;
address_ina = 12;
address_inb = 13;
data_ina = 16'h60;
data_inb = 16'h59;
#10;
address_ina = 14;
address_inb = 15;
data_ina = 16'hfa33;
data_inb = 16'h67b;
#10;
address_ina = 16;
address_inb = 17;
data_ina = 16'hfb8b;
data_inb = 16'hfd38;
#10;
address_ina = 18;
address_inb = 19;
data_ina = 16'hfa82;
data_inb = 16'hff;
#10;
address_ina = 20;
address_inb = 21;
data_ina = 16'h603;
data_inb = 16'h3fa;
#10;
address_ina = 22;
address_inb = 23;
data_ina = 16'hf999;
data_inb = 16'hfc01;
#10;
address_ina = 24;
address_inb = 25;
data_ina = 16'h2f2;
data_inb = 16'h159;
#10;
address_ina = 26;
address_inb = 27;
data_ina = 16'hfd0b;
data_inb = 16'h339;
#10;
address_ina = 28;
address_inb = 29;
data_ina = 16'hfa9e;
data_inb = 16'h505;
#10;
address_ina = 30;
address_inb = 31;
data_ina = 16'hfe7e;
data_inb = 16'hfdcc;
#10;
address_ina = 32;
address_inb = 33;
data_ina = 16'h34a;
data_inb = 16'hfb3f;
#10;
address_ina = 34;
address_inb = 35;
data_ina = 16'hfb6a;
data_inb = 16'h17a;
#10;
address_ina = 36;
address_inb = 37;
data_ina = 16'h33c;
data_inb = 16'h608;
#10;
address_ina = 38;
address_inb = 39;
data_ina = 16'h181;
data_inb = 16'hff88;
#10;
address_ina = 40;
address_inb = 41;
data_ina = 16'hfd7e;
data_inb = 16'hff1e;
#10;
address_ina = 42;
address_inb = 43;
data_ina = 16'h5be;
data_inb = 16'h580;
#10;
address_ina = 44;
address_inb = 45;
data_ina = 16'h66c;
data_inb = 16'hfaed;
#10;
address_ina = 46;
address_inb = 47;
data_ina = 16'h4a1;
data_inb = 16'hfd15;
#10;
address_ina = 48;
address_inb = 49;
data_ina = 16'hfff1;
data_inb = 16'hfb55;
#10;
address_ina = 50;
address_inb = 51;
data_ina = 16'h174;
data_inb = 16'hfc83;
#10;
address_ina = 52;
address_inb = 53;
data_ina = 16'hfe72;
data_inb = 16'hffa9;
#10;
address_ina = 54;
address_inb = 55;
data_ina = 16'hfdab;
data_inb = 16'h5b5;
#10;
address_ina = 56;
address_inb = 57;
data_ina = 16'hfcdd;
data_inb = 16'h1a8;
#10;
address_ina = 58;
address_inb = 59;
data_ina = 16'hfef2;
data_inb = 16'hfd41;
#10;
address_ina = 60;
address_inb = 61;
data_ina = 16'hfd75;
data_inb = 16'hfd52;
#10;
address_ina = 62;
address_inb = 63;
data_ina = 16'hfa16;
data_inb = 16'hfaee;
#10;
address_ina = 64;
address_inb = 65;
data_ina = 16'hff47;
data_inb = 16'h331;
#10;
address_ina = 66;
address_inb = 67;
data_ina = 16'hfe8c;
data_inb = 16'hfea3;
#10;
address_ina = 68;
address_inb = 69;
data_ina = 16'hffa3;
data_inb = 16'hba;
#10;
address_ina = 70;
address_inb = 71;
data_ina = 16'h19;
data_inb = 16'hfad0;
#10;
address_ina = 72;
address_inb = 73;
data_ina = 16'hff5c;
data_inb = 16'h4e4;
#10;
address_ina = 74;
address_inb = 75;
data_ina = 16'h2e;
data_inb = 16'h645;
#10;
address_ina = 76;
address_inb = 77;
data_ina = 16'hfebf;
data_inb = 16'hffaa;
#10;
address_ina = 78;
address_inb = 79;
data_ina = 16'hfee0;
data_inb = 16'h42;
#10;
address_ina = 80;
address_inb = 81;
data_ina = 16'h361;
data_inb = 16'hffec;
#10;
address_ina = 82;
address_inb = 83;
data_ina = 16'hff68;
data_inb = 16'hfb49;
#10;
address_ina = 84;
address_inb = 85;
data_ina = 16'hfa28;
data_inb = 16'h20;
#10;
address_ina = 86;
address_inb = 87;
data_ina = 16'hfdd1;
data_inb = 16'hfc77;
#10;
address_ina = 88;
address_inb = 89;
data_ina = 16'hfdd5;
data_inb = 16'hfd40;
#10;
address_ina = 90;
address_inb = 91;
data_ina = 16'hfa94;
data_inb = 16'hfaab;
#10;
address_ina = 92;
address_inb = 93;
data_ina = 16'hf9a1;
data_inb = 16'hff9c;
#10;
address_ina = 94;
address_inb = 95;
data_ina = 16'h2f9;
data_inb = 16'hfc77;
#10;
address_ina = 96;
address_inb = 97;
data_ina = 16'hfc13;
data_inb = 16'h442;
#10;
address_ina = 98;
address_inb = 99;
data_ina = 16'hfbc9;
data_inb = 16'hfbcf;
#10;
address_ina = 100;
address_inb = 101;
data_ina = 16'h13f;
data_inb = 16'hfc34;
#10;
address_ina = 102;
address_inb = 103;
data_ina = 16'h1ed;
data_inb = 16'h104;
#10;
address_ina = 104;
address_inb = 105;
data_ina = 16'h1c2;
data_inb = 16'hfad7;
#10;
address_ina = 106;
address_inb = 107;
data_ina = 16'hfbb2;
data_inb = 16'hfc38;
#10;
address_ina = 108;
address_inb = 109;
data_ina = 16'hfe33;
data_inb = 16'hfb40;
#10;
address_ina = 110;
address_inb = 111;
data_ina = 16'hfaba;
data_inb = 16'h12;
#10;
address_ina = 112;
address_inb = 113;
data_ina = 16'hf98b;
data_inb = 16'h44c;
#10;
address_ina = 114;
address_inb = 115;
data_ina = 16'h310;
data_inb = 16'hff4e;
#10;
address_ina = 116;
address_inb = 117;
data_ina = 16'hfb5a;
data_inb = 16'h32e;
#10;
address_ina = 118;
address_inb = 119;
data_ina = 16'hfb6f;
data_inb = 16'hfbf1;
#10;
address_ina = 120;
address_inb = 121;
data_ina = 16'hff4c;
data_inb = 16'hfe0d;
#10;
address_ina = 122;
address_inb = 123;
data_ina = 16'hfe0a;
data_inb = 16'hfdd3;
#10;
address_ina = 124;
address_inb = 125;
data_ina = 16'hfaaa;
data_inb = 16'hfe15;
#10;
address_ina = 126;
address_inb = 127;
data_ina = 16'h412;
data_inb = 16'hfc2f;
#10;
address_ina = 128;
address_inb = 129;
data_ina = 16'hfa41;
data_inb = 16'hf9cd;
#10;
address_ina = 130;
address_inb = 131;
data_ina = 16'h32a;
data_inb = 16'h5e5;
#10;
address_ina = 132;
address_inb = 133;
data_ina = 16'h297;
data_inb = 16'h1a2;
#10;
address_ina = 134;
address_inb = 135;
data_ina = 16'hfb90;
data_inb = 16'h60f;
#10;
address_ina = 136;
address_inb = 137;
data_ina = 16'hfecb;
data_inb = 16'h27b;
#10;
address_ina = 138;
address_inb = 139;
data_ina = 16'hfaf2;
data_inb = 16'h310;
#10;
address_ina = 140;
address_inb = 141;
data_ina = 16'h390;
data_inb = 16'hfe6d;
#10;
address_ina = 142;
address_inb = 143;
data_ina = 16'h4cf;
data_inb = 16'h427;
#10;
address_ina = 144;
address_inb = 145;
data_ina = 16'hf9e2;
data_inb = 16'h134;
#10;
address_ina = 146;
address_inb = 147;
data_ina = 16'hfc28;
data_inb = 16'h565;
#10;
address_ina = 148;
address_inb = 149;
data_ina = 16'hfacd;
data_inb = 16'hfc70;
#10;
address_ina = 150;
address_inb = 151;
data_ina = 16'h3c2;
data_inb = 16'hfd7e;
#10;
address_ina = 152;
address_inb = 153;
data_ina = 16'hfd32;
data_inb = 16'hf9f7;
#10;
address_ina = 154;
address_inb = 155;
data_ina = 16'h560;
data_inb = 16'hf9ab;
#10;
address_ina = 156;
address_inb = 157;
data_ina = 16'hfabe;
data_inb = 16'h5b7;
#10;
address_ina = 158;
address_inb = 159;
data_ina = 16'hfd2b;
data_inb = 16'hfe93;
#10;
address_ina = 160;
address_inb = 161;
data_ina = 16'h49;
data_inb = 16'h2d3;
#10;
address_ina = 162;
address_inb = 163;
data_ina = 16'h51a;
data_inb = 16'h348;
#10;
address_ina = 164;
address_inb = 165;
data_ina = 16'h23f;
data_inb = 16'h3cb;
#10;
address_ina = 166;
address_inb = 167;
data_ina = 16'hfb27;
data_inb = 16'hff08;
#10;
address_ina = 168;
address_inb = 169;
data_ina = 16'hfb41;
data_inb = 16'hfd0e;
#10;
address_ina = 170;
address_inb = 171;
data_ina = 16'hff7f;
data_inb = 16'h661;
#10;
address_ina = 172;
address_inb = 173;
data_ina = 16'had;
data_inb = 16'h54;
#10;
address_ina = 174;
address_inb = 175;
data_ina = 16'hfffd;
data_inb = 16'hfb61;
#10;
address_ina = 176;
address_inb = 177;
data_ina = 16'hfd29;
data_inb = 16'hfabb;
#10;
address_ina = 178;
address_inb = 179;
data_ina = 16'hd8;
data_inb = 16'hfeff;
#10;
address_ina = 180;
address_inb = 181;
data_ina = 16'h445;
data_inb = 16'hfddb;
#10;
address_ina = 182;
address_inb = 183;
data_ina = 16'he3;
data_inb = 16'h520;
#10;
address_ina = 184;
address_inb = 185;
data_ina = 16'hfc35;
data_inb = 16'hff26;
#10;
address_ina = 186;
address_inb = 187;
data_ina = 16'hfab5;
data_inb = 16'h208;
#10;
address_ina = 188;
address_inb = 189;
data_ina = 16'hfe3d;
data_inb = 16'h191;
#10;
address_ina = 190;
address_inb = 191;
data_ina = 16'hfbb2;
data_inb = 16'hfab5;
#10;
address_ina = 192;
address_inb = 193;
data_ina = 16'hfa85;
data_inb = 16'h494;
#10;
address_ina = 194;
address_inb = 195;
data_ina = 16'hfb7a;
data_inb = 16'h463;
#10;
address_ina = 196;
address_inb = 197;
data_ina = 16'hfb6b;
data_inb = 16'h101;
#10;
address_ina = 198;
address_inb = 199;
data_ina = 16'h15d;
data_inb = 16'h593;
#10;
address_ina = 200;
address_inb = 201;
data_ina = 16'h29e;
data_inb = 16'hfa67;
#10;
address_ina = 202;
address_inb = 203;
data_ina = 16'h25d;
data_inb = 16'hfd87;
#10;
address_ina = 204;
address_inb = 205;
data_ina = 16'hef;
data_inb = 16'h373;
#10;
address_ina = 206;
address_inb = 207;
data_ina = 16'h210;
data_inb = 16'h5da;
#10;
address_ina = 208;
address_inb = 209;
data_ina = 16'hfd8b;
data_inb = 16'hff8d;
#10;
address_ina = 210;
address_inb = 211;
data_ina = 16'hf985;
data_inb = 16'hfa38;
#10;
address_ina = 212;
address_inb = 213;
data_ina = 16'h1e4;
data_inb = 16'h65a;
#10;
address_ina = 214;
address_inb = 215;
data_ina = 16'hfa19;
data_inb = 16'h23d;
#10;
address_ina = 216;
address_inb = 217;
data_ina = 16'h249;
data_inb = 16'hfcd4;
#10;
address_ina = 218;
address_inb = 219;
data_ina = 16'hfc8d;
data_inb = 16'hfa0f;
#10;
address_ina = 220;
address_inb = 221;
data_ina = 16'h537;
data_inb = 16'hfa46;
#10;
address_ina = 222;
address_inb = 223;
data_ina = 16'hfd49;
data_inb = 16'hfecb;
#10;
address_ina = 224;
address_inb = 225;
data_ina = 16'h5c2;
data_inb = 16'hfe4a;
#10;
address_ina = 226;
address_inb = 227;
data_ina = 16'h174;
data_inb = 16'hfb0e;
#10;
address_ina = 228;
address_inb = 229;
data_ina = 16'h410;
data_inb = 16'hfe16;
#10;
address_ina = 230;
address_inb = 231;
data_ina = 16'h0;
data_inb = 16'h478;
#10;
address_ina = 232;
address_inb = 233;
data_ina = 16'h1bc;
data_inb = 16'h57d;
#10;
address_ina = 234;
address_inb = 235;
data_ina = 16'h3cc;
data_inb = 16'h275;
#10;
address_ina = 236;
address_inb = 237;
data_ina = 16'hfd2d;
data_inb = 16'hfd60;
#10;
address_ina = 238;
address_inb = 239;
data_ina = 16'h1dc;
data_inb = 16'h36c;
#10;
address_ina = 240;
address_inb = 241;
data_ina = 16'hfac3;
data_inb = 16'h132;
#10;
address_ina = 242;
address_inb = 243;
data_ina = 16'h568;
data_inb = 16'h67;
#10;
address_ina = 244;
address_inb = 245;
data_ina = 16'h3de;
data_inb = 16'hfc10;
#10;
address_ina = 246;
address_inb = 247;
data_ina = 16'h156;
data_inb = 16'h4a5;
#10;
address_ina = 248;
address_inb = 249;
data_ina = 16'hfe84;
data_inb = 16'h5c1;
#10;
address_ina = 250;
address_inb = 251;
data_ina = 16'hfab5;
data_inb = 16'h53d;
#10;
address_ina = 252;
address_inb = 253;
data_ina = 16'hfc4b;
data_inb = 16'hfd07;
#10;
address_ina = 254;
address_inb = 255;
data_ina = 16'hfb6a;
data_inb = 16'h15d;
#10;
        wait(init_done);
        #30
        we = 0;
        // Start processing
         
		  #38000

        start = 0;



//        wait (wr_req);
//		  wait (!wr_req);
//		   rd_req = 1;
		  wait(done);
		  #20000
rd_req = 1;
        #70 
		  start = 1;
		 #80 
wait(rd_empty)
rd_req = 0;

$display("Finished the NTT test Number %d",test_num);
////Begin test number #17//////////////
rst = 1;

//#1000
start = 1;
mode = 0; //NTT 0 // INTT 1

// Reset for a few clock cycles

#1000

rst = 0;
test_num = test_num + 1;
#1000
we = 1;
address_ina = 0;
address_inb = 1;
data_ina = 16'h2;
data_inb = 16'hfffe;
#10;
address_ina = 2;
address_inb = 3;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 4;
address_inb = 5;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 6;
address_inb = 7;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 8;
address_inb = 9;
data_ina = 16'h3;
data_inb = 16'h0;
#10;
address_ina = 10;
address_inb = 11;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 12;
address_inb = 13;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 14;
address_inb = 15;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 16;
address_inb = 17;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 18;
address_inb = 19;
data_ina = 16'h2;
data_inb = 16'h0;
#10;
address_ina = 20;
address_inb = 21;
data_ina = 16'h0;
data_inb = 16'h2;
#10;
address_ina = 22;
address_inb = 23;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 24;
address_inb = 25;
data_ina = 16'h2;
data_inb = 16'hfffe;
#10;
address_ina = 26;
address_inb = 27;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 28;
address_inb = 29;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 30;
address_inb = 31;
data_ina = 16'hfffe;
data_inb = 16'hffff;
#10;
address_ina = 32;
address_inb = 33;
data_ina = 16'h0;
data_inb = 16'hfffe;
#10;
address_ina = 34;
address_inb = 35;
data_ina = 16'hfffe;
data_inb = 16'hffff;
#10;
address_ina = 36;
address_inb = 37;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 38;
address_inb = 39;
data_ina = 16'hfffe;
data_inb = 16'h0;
#10;
address_ina = 40;
address_inb = 41;
data_ina = 16'hfffe;
data_inb = 16'h1;
#10;
address_ina = 42;
address_inb = 43;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 44;
address_inb = 45;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 46;
address_inb = 47;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 48;
address_inb = 49;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 50;
address_inb = 51;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 52;
address_inb = 53;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 54;
address_inb = 55;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 56;
address_inb = 57;
data_ina = 16'hfffe;
data_inb = 16'h1;
#10;
address_ina = 58;
address_inb = 59;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 60;
address_inb = 61;
data_ina = 16'h1;
data_inb = 16'h2;
#10;
address_ina = 62;
address_inb = 63;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 64;
address_inb = 65;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 66;
address_inb = 67;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 68;
address_inb = 69;
data_ina = 16'h2;
data_inb = 16'h0;
#10;
address_ina = 70;
address_inb = 71;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 72;
address_inb = 73;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 74;
address_inb = 75;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 76;
address_inb = 77;
data_ina = 16'hfffe;
data_inb = 16'h0;
#10;
address_ina = 78;
address_inb = 79;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 80;
address_inb = 81;
data_ina = 16'h2;
data_inb = 16'h1;
#10;
address_ina = 82;
address_inb = 83;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 84;
address_inb = 85;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 86;
address_inb = 87;
data_ina = 16'h2;
data_inb = 16'hfffe;
#10;
address_ina = 88;
address_inb = 89;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 90;
address_inb = 91;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 92;
address_inb = 93;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 94;
address_inb = 95;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 96;
address_inb = 97;
data_ina = 16'h2;
data_inb = 16'h1;
#10;
address_ina = 98;
address_inb = 99;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 100;
address_inb = 101;
data_ina = 16'h0;
data_inb = 16'h2;
#10;
address_ina = 102;
address_inb = 103;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 104;
address_inb = 105;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 106;
address_inb = 107;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 108;
address_inb = 109;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 110;
address_inb = 111;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 112;
address_inb = 113;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 114;
address_inb = 115;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 116;
address_inb = 117;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 118;
address_inb = 119;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 120;
address_inb = 121;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 122;
address_inb = 123;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 124;
address_inb = 125;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 126;
address_inb = 127;
data_ina = 16'hffff;
data_inb = 16'h2;
#10;
address_ina = 128;
address_inb = 129;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 130;
address_inb = 131;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 132;
address_inb = 133;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 134;
address_inb = 135;
data_ina = 16'h2;
data_inb = 16'h1;
#10;
address_ina = 136;
address_inb = 137;
data_ina = 16'hfffe;
data_inb = 16'h0;
#10;
address_ina = 138;
address_inb = 139;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 140;
address_inb = 141;
data_ina = 16'h1;
data_inb = 16'hfffd;
#10;
address_ina = 142;
address_inb = 143;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 144;
address_inb = 145;
data_ina = 16'hfffe;
data_inb = 16'hffff;
#10;
address_ina = 146;
address_inb = 147;
data_ina = 16'h2;
data_inb = 16'h2;
#10;
address_ina = 148;
address_inb = 149;
data_ina = 16'hfffd;
data_inb = 16'hffff;
#10;
address_ina = 150;
address_inb = 151;
data_ina = 16'hfffe;
data_inb = 16'hfffe;
#10;
address_ina = 152;
address_inb = 153;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 154;
address_inb = 155;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 156;
address_inb = 157;
data_ina = 16'hfffe;
data_inb = 16'h1;
#10;
address_ina = 158;
address_inb = 159;
data_ina = 16'h2;
data_inb = 16'h0;
#10;
address_ina = 160;
address_inb = 161;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 162;
address_inb = 163;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 164;
address_inb = 165;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 166;
address_inb = 167;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 168;
address_inb = 169;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 170;
address_inb = 171;
data_ina = 16'hfffe;
data_inb = 16'hffff;
#10;
address_ina = 172;
address_inb = 173;
data_ina = 16'h1;
data_inb = 16'hfffe;
#10;
address_ina = 174;
address_inb = 175;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 176;
address_inb = 177;
data_ina = 16'hfffe;
data_inb = 16'hfffe;
#10;
address_ina = 178;
address_inb = 179;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 180;
address_inb = 181;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 182;
address_inb = 183;
data_ina = 16'hfffe;
data_inb = 16'h0;
#10;
address_ina = 184;
address_inb = 185;
data_ina = 16'h0;
data_inb = 16'hfffe;
#10;
address_ina = 186;
address_inb = 187;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 188;
address_inb = 189;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 190;
address_inb = 191;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 192;
address_inb = 193;
data_ina = 16'hfffd;
data_inb = 16'h1;
#10;
address_ina = 194;
address_inb = 195;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 196;
address_inb = 197;
data_ina = 16'h1;
data_inb = 16'h2;
#10;
address_ina = 198;
address_inb = 199;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 200;
address_inb = 201;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 202;
address_inb = 203;
data_ina = 16'hfffe;
data_inb = 16'h1;
#10;
address_ina = 204;
address_inb = 205;
data_ina = 16'hffff;
data_inb = 16'hfffe;
#10;
address_ina = 206;
address_inb = 207;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 208;
address_inb = 209;
data_ina = 16'h2;
data_inb = 16'h0;
#10;
address_ina = 210;
address_inb = 211;
data_ina = 16'hfffe;
data_inb = 16'h1;
#10;
address_ina = 212;
address_inb = 213;
data_ina = 16'hffff;
data_inb = 16'hfffe;
#10;
address_ina = 214;
address_inb = 215;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 216;
address_inb = 217;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 218;
address_inb = 219;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 220;
address_inb = 221;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 222;
address_inb = 223;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 224;
address_inb = 225;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 226;
address_inb = 227;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 228;
address_inb = 229;
data_ina = 16'h2;
data_inb = 16'h2;
#10;
address_ina = 230;
address_inb = 231;
data_ina = 16'h2;
data_inb = 16'hfffe;
#10;
address_ina = 232;
address_inb = 233;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 234;
address_inb = 235;
data_ina = 16'h1;
data_inb = 16'hfffe;
#10;
address_ina = 236;
address_inb = 237;
data_ina = 16'h2;
data_inb = 16'hffff;
#10;
address_ina = 238;
address_inb = 239;
data_ina = 16'h3;
data_inb = 16'hffff;
#10;
address_ina = 240;
address_inb = 241;
data_ina = 16'hfffe;
data_inb = 16'hffff;
#10;
address_ina = 242;
address_inb = 243;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 244;
address_inb = 245;
data_ina = 16'h0;
data_inb = 16'h2;
#10;
address_ina = 246;
address_inb = 247;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 248;
address_inb = 249;
data_ina = 16'hfffe;
data_inb = 16'h1;
#10;
address_ina = 250;
address_inb = 251;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 252;
address_inb = 253;
data_ina = 16'hfffe;
data_inb = 16'hfffe;
#10;
address_ina = 254;
address_inb = 255;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
        wait(init_done);
        #30
        we = 0;
        // Start processing
         
		  #38000

        start = 0;



//        wait (wr_req);
//		  wait (!wr_req);
//		   rd_req = 1;
		  wait(done);
		  #20000
rd_req = 1;
        #70 
		  start = 1;
		 #80 
wait(rd_empty)
rd_req = 0;

$display("Finished the NTT test Number %d",test_num);
////Begin test number #18//////////////
rst = 1;

//#1000
start = 1;
mode = 0; //NTT 0 // INTT 1

// Reset for a few clock cycles

#1000

rst = 0;
test_num = test_num + 1;
#1000
we = 1;
address_ina = 0;
address_inb = 1;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 2;
address_inb = 3;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 4;
address_inb = 5;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 6;
address_inb = 7;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 8;
address_inb = 9;
data_ina = 16'h2;
data_inb = 16'h2;
#10;
address_ina = 10;
address_inb = 11;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 12;
address_inb = 13;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 14;
address_inb = 15;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 16;
address_inb = 17;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 18;
address_inb = 19;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 20;
address_inb = 21;
data_ina = 16'h2;
data_inb = 16'h0;
#10;
address_ina = 22;
address_inb = 23;
data_ina = 16'h2;
data_inb = 16'h2;
#10;
address_ina = 24;
address_inb = 25;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 26;
address_inb = 27;
data_ina = 16'hfffe;
data_inb = 16'h0;
#10;
address_ina = 28;
address_inb = 29;
data_ina = 16'hfffe;
data_inb = 16'h3;
#10;
address_ina = 30;
address_inb = 31;
data_ina = 16'h2;
data_inb = 16'h1;
#10;
address_ina = 32;
address_inb = 33;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 34;
address_inb = 35;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 36;
address_inb = 37;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 38;
address_inb = 39;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 40;
address_inb = 41;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 42;
address_inb = 43;
data_ina = 16'h2;
data_inb = 16'h1;
#10;
address_ina = 44;
address_inb = 45;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 46;
address_inb = 47;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 48;
address_inb = 49;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 50;
address_inb = 51;
data_ina = 16'h2;
data_inb = 16'h2;
#10;
address_ina = 52;
address_inb = 53;
data_ina = 16'hfffe;
data_inb = 16'h2;
#10;
address_ina = 54;
address_inb = 55;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 56;
address_inb = 57;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 58;
address_inb = 59;
data_ina = 16'h0;
data_inb = 16'h2;
#10;
address_ina = 60;
address_inb = 61;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 62;
address_inb = 63;
data_ina = 16'hfffe;
data_inb = 16'hffff;
#10;
address_ina = 64;
address_inb = 65;
data_ina = 16'hffff;
data_inb = 16'hfffe;
#10;
address_ina = 66;
address_inb = 67;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 68;
address_inb = 69;
data_ina = 16'hfffe;
data_inb = 16'h0;
#10;
address_ina = 70;
address_inb = 71;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 72;
address_inb = 73;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 74;
address_inb = 75;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 76;
address_inb = 77;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 78;
address_inb = 79;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 80;
address_inb = 81;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 82;
address_inb = 83;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 84;
address_inb = 85;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 86;
address_inb = 87;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 88;
address_inb = 89;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 90;
address_inb = 91;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 92;
address_inb = 93;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 94;
address_inb = 95;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 96;
address_inb = 97;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 98;
address_inb = 99;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 100;
address_inb = 101;
data_ina = 16'h1;
data_inb = 16'h2;
#10;
address_ina = 102;
address_inb = 103;
data_ina = 16'hfffe;
data_inb = 16'hffff;
#10;
address_ina = 104;
address_inb = 105;
data_ina = 16'hfffe;
data_inb = 16'h0;
#10;
address_ina = 106;
address_inb = 107;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 108;
address_inb = 109;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 110;
address_inb = 111;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 112;
address_inb = 113;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 114;
address_inb = 115;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 116;
address_inb = 117;
data_ina = 16'h2;
data_inb = 16'hffff;
#10;
address_ina = 118;
address_inb = 119;
data_ina = 16'h2;
data_inb = 16'h2;
#10;
address_ina = 120;
address_inb = 121;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 122;
address_inb = 123;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 124;
address_inb = 125;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 126;
address_inb = 127;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 128;
address_inb = 129;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 130;
address_inb = 131;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 132;
address_inb = 133;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 134;
address_inb = 135;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 136;
address_inb = 137;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 138;
address_inb = 139;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 140;
address_inb = 141;
data_ina = 16'h3;
data_inb = 16'h2;
#10;
address_ina = 142;
address_inb = 143;
data_ina = 16'h2;
data_inb = 16'h1;
#10;
address_ina = 144;
address_inb = 145;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 146;
address_inb = 147;
data_ina = 16'hffff;
data_inb = 16'hfffe;
#10;
address_ina = 148;
address_inb = 149;
data_ina = 16'hfffd;
data_inb = 16'h1;
#10;
address_ina = 150;
address_inb = 151;
data_ina = 16'h0;
data_inb = 16'h2;
#10;
address_ina = 152;
address_inb = 153;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 154;
address_inb = 155;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 156;
address_inb = 157;
data_ina = 16'h0;
data_inb = 16'hfffe;
#10;
address_ina = 158;
address_inb = 159;
data_ina = 16'h0;
data_inb = 16'h2;
#10;
address_ina = 160;
address_inb = 161;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 162;
address_inb = 163;
data_ina = 16'hfffe;
data_inb = 16'h0;
#10;
address_ina = 164;
address_inb = 165;
data_ina = 16'hfffe;
data_inb = 16'h1;
#10;
address_ina = 166;
address_inb = 167;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 168;
address_inb = 169;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 170;
address_inb = 171;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 172;
address_inb = 173;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 174;
address_inb = 175;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 176;
address_inb = 177;
data_ina = 16'h1;
data_inb = 16'hfffe;
#10;
address_ina = 178;
address_inb = 179;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 180;
address_inb = 181;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 182;
address_inb = 183;
data_ina = 16'h2;
data_inb = 16'h1;
#10;
address_ina = 184;
address_inb = 185;
data_ina = 16'hfffe;
data_inb = 16'hfffe;
#10;
address_ina = 186;
address_inb = 187;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 188;
address_inb = 189;
data_ina = 16'h1;
data_inb = 16'hfffe;
#10;
address_ina = 190;
address_inb = 191;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 192;
address_inb = 193;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 194;
address_inb = 195;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 196;
address_inb = 197;
data_ina = 16'hffff;
data_inb = 16'h2;
#10;
address_ina = 198;
address_inb = 199;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 200;
address_inb = 201;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 202;
address_inb = 203;
data_ina = 16'hffff;
data_inb = 16'hfffe;
#10;
address_ina = 204;
address_inb = 205;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 206;
address_inb = 207;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 208;
address_inb = 209;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 210;
address_inb = 211;
data_ina = 16'h1;
data_inb = 16'h2;
#10;
address_ina = 212;
address_inb = 213;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 214;
address_inb = 215;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 216;
address_inb = 217;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 218;
address_inb = 219;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 220;
address_inb = 221;
data_ina = 16'hfffd;
data_inb = 16'hffff;
#10;
address_ina = 222;
address_inb = 223;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 224;
address_inb = 225;
data_ina = 16'h2;
data_inb = 16'hffff;
#10;
address_ina = 226;
address_inb = 227;
data_ina = 16'h1;
data_inb = 16'hfffe;
#10;
address_ina = 228;
address_inb = 229;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 230;
address_inb = 231;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 232;
address_inb = 233;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 234;
address_inb = 235;
data_ina = 16'h2;
data_inb = 16'h1;
#10;
address_ina = 236;
address_inb = 237;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 238;
address_inb = 239;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 240;
address_inb = 241;
data_ina = 16'hfffe;
data_inb = 16'h2;
#10;
address_ina = 242;
address_inb = 243;
data_ina = 16'hffff;
data_inb = 16'h2;
#10;
address_ina = 244;
address_inb = 245;
data_ina = 16'h0;
data_inb = 16'hfffe;
#10;
address_ina = 246;
address_inb = 247;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 248;
address_inb = 249;
data_ina = 16'hfffe;
data_inb = 16'h0;
#10;
address_ina = 250;
address_inb = 251;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 252;
address_inb = 253;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 254;
address_inb = 255;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
        wait(init_done);
        #30
        we = 0;
        // Start processing
         
		  #38000

        start = 0;



//        wait (wr_req);
//		  wait (!wr_req);
//		   rd_req = 1;
		  wait(done);
		  #20000
rd_req = 1;
        #70 
		  start = 1;
		 #80 
wait(rd_empty)
rd_req = 0;

$display("Finished the NTT test Number %d",test_num);
////Begin test number #19//////////////
rst = 1;

//#1000
start = 1;
mode = 0; //NTT 0 // INTT 1

// Reset for a few clock cycles

#1000

rst = 0;
test_num = test_num + 1;
#1000
we = 1;
address_ina = 0;
address_inb = 1;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 2;
address_inb = 3;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 4;
address_inb = 5;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 6;
address_inb = 7;
data_ina = 16'h0;
data_inb = 16'hfffd;
#10;
address_ina = 8;
address_inb = 9;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 10;
address_inb = 11;
data_ina = 16'h2;
data_inb = 16'h2;
#10;
address_ina = 12;
address_inb = 13;
data_ina = 16'h0;
data_inb = 16'hfffe;
#10;
address_ina = 14;
address_inb = 15;
data_ina = 16'hfffe;
data_inb = 16'h0;
#10;
address_ina = 16;
address_inb = 17;
data_ina = 16'hfffe;
data_inb = 16'h1;
#10;
address_ina = 18;
address_inb = 19;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 20;
address_inb = 21;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 22;
address_inb = 23;
data_ina = 16'h0;
data_inb = 16'h2;
#10;
address_ina = 24;
address_inb = 25;
data_ina = 16'h1;
data_inb = 16'hfffe;
#10;
address_ina = 26;
address_inb = 27;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 28;
address_inb = 29;
data_ina = 16'hfffe;
data_inb = 16'h1;
#10;
address_ina = 30;
address_inb = 31;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 32;
address_inb = 33;
data_ina = 16'h1;
data_inb = 16'hfffe;
#10;
address_ina = 34;
address_inb = 35;
data_ina = 16'h0;
data_inb = 16'hfffe;
#10;
address_ina = 36;
address_inb = 37;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 38;
address_inb = 39;
data_ina = 16'h2;
data_inb = 16'hffff;
#10;
address_ina = 40;
address_inb = 41;
data_ina = 16'hfffd;
data_inb = 16'h0;
#10;
address_ina = 42;
address_inb = 43;
data_ina = 16'h0;
data_inb = 16'hfffe;
#10;
address_ina = 44;
address_inb = 45;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 46;
address_inb = 47;
data_ina = 16'h0;
data_inb = 16'h3;
#10;
address_ina = 48;
address_inb = 49;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 50;
address_inb = 51;
data_ina = 16'hfffe;
data_inb = 16'h0;
#10;
address_ina = 52;
address_inb = 53;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 54;
address_inb = 55;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 56;
address_inb = 57;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 58;
address_inb = 59;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 60;
address_inb = 61;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 62;
address_inb = 63;
data_ina = 16'h2;
data_inb = 16'hffff;
#10;
address_ina = 64;
address_inb = 65;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 66;
address_inb = 67;
data_ina = 16'h0;
data_inb = 16'hfffe;
#10;
address_ina = 68;
address_inb = 69;
data_ina = 16'h1;
data_inb = 16'h2;
#10;
address_ina = 70;
address_inb = 71;
data_ina = 16'h0;
data_inb = 16'hfffe;
#10;
address_ina = 72;
address_inb = 73;
data_ina = 16'h2;
data_inb = 16'hfffe;
#10;
address_ina = 74;
address_inb = 75;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 76;
address_inb = 77;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 78;
address_inb = 79;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 80;
address_inb = 81;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 82;
address_inb = 83;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 84;
address_inb = 85;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 86;
address_inb = 87;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 88;
address_inb = 89;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 90;
address_inb = 91;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 92;
address_inb = 93;
data_ina = 16'h2;
data_inb = 16'h1;
#10;
address_ina = 94;
address_inb = 95;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 96;
address_inb = 97;
data_ina = 16'hffff;
data_inb = 16'h3;
#10;
address_ina = 98;
address_inb = 99;
data_ina = 16'hfffe;
data_inb = 16'h0;
#10;
address_ina = 100;
address_inb = 101;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 102;
address_inb = 103;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 104;
address_inb = 105;
data_ina = 16'hfffe;
data_inb = 16'h1;
#10;
address_ina = 106;
address_inb = 107;
data_ina = 16'hfffe;
data_inb = 16'h2;
#10;
address_ina = 108;
address_inb = 109;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 110;
address_inb = 111;
data_ina = 16'hfffd;
data_inb = 16'h0;
#10;
address_ina = 112;
address_inb = 113;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 114;
address_inb = 115;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 116;
address_inb = 117;
data_ina = 16'h2;
data_inb = 16'hfffe;
#10;
address_ina = 118;
address_inb = 119;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 120;
address_inb = 121;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 122;
address_inb = 123;
data_ina = 16'h2;
data_inb = 16'h1;
#10;
address_ina = 124;
address_inb = 125;
data_ina = 16'hfffe;
data_inb = 16'hffff;
#10;
address_ina = 126;
address_inb = 127;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 128;
address_inb = 129;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 130;
address_inb = 131;
data_ina = 16'hfffe;
data_inb = 16'h1;
#10;
address_ina = 132;
address_inb = 133;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 134;
address_inb = 135;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 136;
address_inb = 137;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 138;
address_inb = 139;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 140;
address_inb = 141;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 142;
address_inb = 143;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 144;
address_inb = 145;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 146;
address_inb = 147;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 148;
address_inb = 149;
data_ina = 16'hfffe;
data_inb = 16'hfffe;
#10;
address_ina = 150;
address_inb = 151;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 152;
address_inb = 153;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 154;
address_inb = 155;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 156;
address_inb = 157;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 158;
address_inb = 159;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 160;
address_inb = 161;
data_ina = 16'h1;
data_inb = 16'h2;
#10;
address_ina = 162;
address_inb = 163;
data_ina = 16'hfffe;
data_inb = 16'h1;
#10;
address_ina = 164;
address_inb = 165;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 166;
address_inb = 167;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 168;
address_inb = 169;
data_ina = 16'h2;
data_inb = 16'h0;
#10;
address_ina = 170;
address_inb = 171;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 172;
address_inb = 173;
data_ina = 16'hfffe;
data_inb = 16'h0;
#10;
address_ina = 174;
address_inb = 175;
data_ina = 16'hffff;
data_inb = 16'hfffe;
#10;
address_ina = 176;
address_inb = 177;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 178;
address_inb = 179;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 180;
address_inb = 181;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 182;
address_inb = 183;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 184;
address_inb = 185;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 186;
address_inb = 187;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 188;
address_inb = 189;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 190;
address_inb = 191;
data_ina = 16'hfffe;
data_inb = 16'hffff;
#10;
address_ina = 192;
address_inb = 193;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 194;
address_inb = 195;
data_ina = 16'hfffe;
data_inb = 16'h0;
#10;
address_ina = 196;
address_inb = 197;
data_ina = 16'h0;
data_inb = 16'hfffe;
#10;
address_ina = 198;
address_inb = 199;
data_ina = 16'hffff;
data_inb = 16'h2;
#10;
address_ina = 200;
address_inb = 201;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 202;
address_inb = 203;
data_ina = 16'h3;
data_inb = 16'hfffe;
#10;
address_ina = 204;
address_inb = 205;
data_ina = 16'h2;
data_inb = 16'h0;
#10;
address_ina = 206;
address_inb = 207;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 208;
address_inb = 209;
data_ina = 16'h2;
data_inb = 16'hffff;
#10;
address_ina = 210;
address_inb = 211;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 212;
address_inb = 213;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 214;
address_inb = 215;
data_ina = 16'h3;
data_inb = 16'hfffe;
#10;
address_ina = 216;
address_inb = 217;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 218;
address_inb = 219;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 220;
address_inb = 221;
data_ina = 16'h0;
data_inb = 16'hfffe;
#10;
address_ina = 222;
address_inb = 223;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 224;
address_inb = 225;
data_ina = 16'h0;
data_inb = 16'hfffe;
#10;
address_ina = 226;
address_inb = 227;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 228;
address_inb = 229;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 230;
address_inb = 231;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 232;
address_inb = 233;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 234;
address_inb = 235;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 236;
address_inb = 237;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 238;
address_inb = 239;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 240;
address_inb = 241;
data_ina = 16'h0;
data_inb = 16'h3;
#10;
address_ina = 242;
address_inb = 243;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 244;
address_inb = 245;
data_ina = 16'h2;
data_inb = 16'h0;
#10;
address_ina = 246;
address_inb = 247;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 248;
address_inb = 249;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 250;
address_inb = 251;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 252;
address_inb = 253;
data_ina = 16'h0;
data_inb = 16'hfffe;
#10;
address_ina = 254;
address_inb = 255;
data_ina = 16'h1;
data_inb = 16'h3;
#10;
        wait(init_done);
        #30
        we = 0;
        // Start processing
         
		  #38000

        start = 0;



//        wait (wr_req);
//		  wait (!wr_req);
//		   rd_req = 1;
		  wait(done);
		  #20000
rd_req = 1;
        #70 
		  start = 1;
		 #80 
wait(rd_empty)
rd_req = 0;

$display("Finished the NTT test Number %d",test_num);
////Begin test number #20//////////////
rst = 1;

//#1000
start = 1;
mode = 0; //NTT 0 // INTT 1

// Reset for a few clock cycles

#1000

rst = 0;
test_num = test_num + 1;
#1000
we = 1;
address_ina = 0;
address_inb = 1;
data_ina = 16'hffff;
data_inb = 16'h2;
#10;
address_ina = 2;
address_inb = 3;
data_ina = 16'h2;
data_inb = 16'h0;
#10;
address_ina = 4;
address_inb = 5;
data_ina = 16'h0;
data_inb = 16'h2;
#10;
address_ina = 6;
address_inb = 7;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 8;
address_inb = 9;
data_ina = 16'hfffe;
data_inb = 16'hffff;
#10;
address_ina = 10;
address_inb = 11;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 12;
address_inb = 13;
data_ina = 16'h2;
data_inb = 16'h0;
#10;
address_ina = 14;
address_inb = 15;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 16;
address_inb = 17;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 18;
address_inb = 19;
data_ina = 16'h2;
data_inb = 16'h2;
#10;
address_ina = 20;
address_inb = 21;
data_ina = 16'h0;
data_inb = 16'h2;
#10;
address_ina = 22;
address_inb = 23;
data_ina = 16'h2;
data_inb = 16'hffff;
#10;
address_ina = 24;
address_inb = 25;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 26;
address_inb = 27;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 28;
address_inb = 29;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 30;
address_inb = 31;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 32;
address_inb = 33;
data_ina = 16'hffff;
data_inb = 16'hfffe;
#10;
address_ina = 34;
address_inb = 35;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 36;
address_inb = 37;
data_ina = 16'h0;
data_inb = 16'hfffe;
#10;
address_ina = 38;
address_inb = 39;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 40;
address_inb = 41;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 42;
address_inb = 43;
data_ina = 16'h2;
data_inb = 16'hffff;
#10;
address_ina = 44;
address_inb = 45;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 46;
address_inb = 47;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 48;
address_inb = 49;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 50;
address_inb = 51;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 52;
address_inb = 53;
data_ina = 16'h2;
data_inb = 16'h1;
#10;
address_ina = 54;
address_inb = 55;
data_ina = 16'hfffe;
data_inb = 16'h0;
#10;
address_ina = 56;
address_inb = 57;
data_ina = 16'hfffe;
data_inb = 16'h1;
#10;
address_ina = 58;
address_inb = 59;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 60;
address_inb = 61;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 62;
address_inb = 63;
data_ina = 16'h0;
data_inb = 16'hfffe;
#10;
address_ina = 64;
address_inb = 65;
data_ina = 16'hffff;
data_inb = 16'hfffe;
#10;
address_ina = 66;
address_inb = 67;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 68;
address_inb = 69;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 70;
address_inb = 71;
data_ina = 16'h2;
data_inb = 16'h0;
#10;
address_ina = 72;
address_inb = 73;
data_ina = 16'hfffe;
data_inb = 16'h0;
#10;
address_ina = 74;
address_inb = 75;
data_ina = 16'h2;
data_inb = 16'h0;
#10;
address_ina = 76;
address_inb = 77;
data_ina = 16'hffff;
data_inb = 16'hfffe;
#10;
address_ina = 78;
address_inb = 79;
data_ina = 16'h3;
data_inb = 16'h0;
#10;
address_ina = 80;
address_inb = 81;
data_ina = 16'hfffe;
data_inb = 16'hffff;
#10;
address_ina = 82;
address_inb = 83;
data_ina = 16'h2;
data_inb = 16'hffff;
#10;
address_ina = 84;
address_inb = 85;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 86;
address_inb = 87;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 88;
address_inb = 89;
data_ina = 16'h0;
data_inb = 16'h2;
#10;
address_ina = 90;
address_inb = 91;
data_ina = 16'h2;
data_inb = 16'h0;
#10;
address_ina = 92;
address_inb = 93;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 94;
address_inb = 95;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 96;
address_inb = 97;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 98;
address_inb = 99;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 100;
address_inb = 101;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 102;
address_inb = 103;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 104;
address_inb = 105;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 106;
address_inb = 107;
data_ina = 16'hffff;
data_inb = 16'h2;
#10;
address_ina = 108;
address_inb = 109;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 110;
address_inb = 111;
data_ina = 16'hfffe;
data_inb = 16'h0;
#10;
address_ina = 112;
address_inb = 113;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 114;
address_inb = 115;
data_ina = 16'h0;
data_inb = 16'hfffe;
#10;
address_ina = 116;
address_inb = 117;
data_ina = 16'h0;
data_inb = 16'hfffe;
#10;
address_ina = 118;
address_inb = 119;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 120;
address_inb = 121;
data_ina = 16'h2;
data_inb = 16'h3;
#10;
address_ina = 122;
address_inb = 123;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 124;
address_inb = 125;
data_ina = 16'hffff;
data_inb = 16'h2;
#10;
address_ina = 126;
address_inb = 127;
data_ina = 16'h2;
data_inb = 16'h1;
#10;
address_ina = 128;
address_inb = 129;
data_ina = 16'h0;
data_inb = 16'hfffe;
#10;
address_ina = 130;
address_inb = 131;
data_ina = 16'h2;
data_inb = 16'h0;
#10;
address_ina = 132;
address_inb = 133;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 134;
address_inb = 135;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 136;
address_inb = 137;
data_ina = 16'h1;
data_inb = 16'hfffe;
#10;
address_ina = 138;
address_inb = 139;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 140;
address_inb = 141;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 142;
address_inb = 143;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 144;
address_inb = 145;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 146;
address_inb = 147;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 148;
address_inb = 149;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 150;
address_inb = 151;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 152;
address_inb = 153;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 154;
address_inb = 155;
data_ina = 16'hffff;
data_inb = 16'hfffe;
#10;
address_ina = 156;
address_inb = 157;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 158;
address_inb = 159;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 160;
address_inb = 161;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 162;
address_inb = 163;
data_ina = 16'hfffe;
data_inb = 16'hfffe;
#10;
address_ina = 164;
address_inb = 165;
data_ina = 16'h0;
data_inb = 16'h2;
#10;
address_ina = 166;
address_inb = 167;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 168;
address_inb = 169;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 170;
address_inb = 171;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 172;
address_inb = 173;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 174;
address_inb = 175;
data_ina = 16'hffff;
data_inb = 16'hfffe;
#10;
address_ina = 176;
address_inb = 177;
data_ina = 16'hfffe;
data_inb = 16'h1;
#10;
address_ina = 178;
address_inb = 179;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 180;
address_inb = 181;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 182;
address_inb = 183;
data_ina = 16'h2;
data_inb = 16'h0;
#10;
address_ina = 184;
address_inb = 185;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 186;
address_inb = 187;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 188;
address_inb = 189;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 190;
address_inb = 191;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 192;
address_inb = 193;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 194;
address_inb = 195;
data_ina = 16'hfffe;
data_inb = 16'h0;
#10;
address_ina = 196;
address_inb = 197;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 198;
address_inb = 199;
data_ina = 16'hfffe;
data_inb = 16'h1;
#10;
address_ina = 200;
address_inb = 201;
data_ina = 16'hfffe;
data_inb = 16'hfffe;
#10;
address_ina = 202;
address_inb = 203;
data_ina = 16'h3;
data_inb = 16'h1;
#10;
address_ina = 204;
address_inb = 205;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 206;
address_inb = 207;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 208;
address_inb = 209;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 210;
address_inb = 211;
data_ina = 16'h0;
data_inb = 16'hfffe;
#10;
address_ina = 212;
address_inb = 213;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 214;
address_inb = 215;
data_ina = 16'hffff;
data_inb = 16'h2;
#10;
address_ina = 216;
address_inb = 217;
data_ina = 16'hffff;
data_inb = 16'h2;
#10;
address_ina = 218;
address_inb = 219;
data_ina = 16'h1;
data_inb = 16'h2;
#10;
address_ina = 220;
address_inb = 221;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 222;
address_inb = 223;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 224;
address_inb = 225;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 226;
address_inb = 227;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 228;
address_inb = 229;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 230;
address_inb = 231;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 232;
address_inb = 233;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 234;
address_inb = 235;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 236;
address_inb = 237;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 238;
address_inb = 239;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 240;
address_inb = 241;
data_ina = 16'h2;
data_inb = 16'hffff;
#10;
address_ina = 242;
address_inb = 243;
data_ina = 16'hffff;
data_inb = 16'hfffe;
#10;
address_ina = 244;
address_inb = 245;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 246;
address_inb = 247;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 248;
address_inb = 249;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 250;
address_inb = 251;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 252;
address_inb = 253;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 254;
address_inb = 255;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
        wait(init_done);
        #30
        we = 0;
        // Start processing
         
		  #38000

        start = 0;



//        wait (wr_req);
//		  wait (!wr_req);
//		   rd_req = 1;
		  wait(done);
		  #20000
rd_req = 1;
        #70 
		  start = 1;
		 #80 
wait(rd_empty)
rd_req = 0;

$display("Finished the NTT test Number %d",test_num);
////Begin test number #21//////////////
rst = 1;

//#1000
start = 1;
mode = 0; //NTT 0 // INTT 1

// Reset for a few clock cycles

#1000

rst = 0;
test_num = test_num + 1;
#1000
we = 1;
address_ina = 0;
address_inb = 1;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 2;
address_inb = 3;
data_ina = 16'h2;
data_inb = 16'h0;
#10;
address_ina = 4;
address_inb = 5;
data_ina = 16'h1;
data_inb = 16'h2;
#10;
address_ina = 6;
address_inb = 7;
data_ina = 16'hfffe;
data_inb = 16'h0;
#10;
address_ina = 8;
address_inb = 9;
data_ina = 16'h2;
data_inb = 16'h1;
#10;
address_ina = 10;
address_inb = 11;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 12;
address_inb = 13;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 14;
address_inb = 15;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 16;
address_inb = 17;
data_ina = 16'h1;
data_inb = 16'h2;
#10;
address_ina = 18;
address_inb = 19;
data_ina = 16'h1;
data_inb = 16'hfffe;
#10;
address_ina = 20;
address_inb = 21;
data_ina = 16'hfffe;
data_inb = 16'hffff;
#10;
address_ina = 22;
address_inb = 23;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 24;
address_inb = 25;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 26;
address_inb = 27;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 28;
address_inb = 29;
data_ina = 16'hfffe;
data_inb = 16'h1;
#10;
address_ina = 30;
address_inb = 31;
data_ina = 16'h0;
data_inb = 16'h2;
#10;
address_ina = 32;
address_inb = 33;
data_ina = 16'h2;
data_inb = 16'h1;
#10;
address_ina = 34;
address_inb = 35;
data_ina = 16'hffff;
data_inb = 16'hfffe;
#10;
address_ina = 36;
address_inb = 37;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 38;
address_inb = 39;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 40;
address_inb = 41;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 42;
address_inb = 43;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 44;
address_inb = 45;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 46;
address_inb = 47;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 48;
address_inb = 49;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 50;
address_inb = 51;
data_ina = 16'hffff;
data_inb = 16'hfffe;
#10;
address_ina = 52;
address_inb = 53;
data_ina = 16'hfffe;
data_inb = 16'h0;
#10;
address_ina = 54;
address_inb = 55;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 56;
address_inb = 57;
data_ina = 16'h0;
data_inb = 16'h2;
#10;
address_ina = 58;
address_inb = 59;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 60;
address_inb = 61;
data_ina = 16'hfffe;
data_inb = 16'hffff;
#10;
address_ina = 62;
address_inb = 63;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 64;
address_inb = 65;
data_ina = 16'h3;
data_inb = 16'hfffe;
#10;
address_ina = 66;
address_inb = 67;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 68;
address_inb = 69;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 70;
address_inb = 71;
data_ina = 16'h0;
data_inb = 16'h3;
#10;
address_ina = 72;
address_inb = 73;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 74;
address_inb = 75;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 76;
address_inb = 77;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 78;
address_inb = 79;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 80;
address_inb = 81;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 82;
address_inb = 83;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 84;
address_inb = 85;
data_ina = 16'h2;
data_inb = 16'h0;
#10;
address_ina = 86;
address_inb = 87;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 88;
address_inb = 89;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 90;
address_inb = 91;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 92;
address_inb = 93;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 94;
address_inb = 95;
data_ina = 16'hfffe;
data_inb = 16'h0;
#10;
address_ina = 96;
address_inb = 97;
data_ina = 16'hfffe;
data_inb = 16'h0;
#10;
address_ina = 98;
address_inb = 99;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 100;
address_inb = 101;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 102;
address_inb = 103;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 104;
address_inb = 105;
data_ina = 16'h2;
data_inb = 16'h0;
#10;
address_ina = 106;
address_inb = 107;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 108;
address_inb = 109;
data_ina = 16'h1;
data_inb = 16'hfffe;
#10;
address_ina = 110;
address_inb = 111;
data_ina = 16'h2;
data_inb = 16'hffff;
#10;
address_ina = 112;
address_inb = 113;
data_ina = 16'hfffe;
data_inb = 16'hfffe;
#10;
address_ina = 114;
address_inb = 115;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 116;
address_inb = 117;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 118;
address_inb = 119;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 120;
address_inb = 121;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 122;
address_inb = 123;
data_ina = 16'hfffd;
data_inb = 16'hffff;
#10;
address_ina = 124;
address_inb = 125;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 126;
address_inb = 127;
data_ina = 16'hffff;
data_inb = 16'h2;
#10;
address_ina = 128;
address_inb = 129;
data_ina = 16'hfffe;
data_inb = 16'h2;
#10;
address_ina = 130;
address_inb = 131;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 132;
address_inb = 133;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 134;
address_inb = 135;
data_ina = 16'hfffe;
data_inb = 16'hffff;
#10;
address_ina = 136;
address_inb = 137;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 138;
address_inb = 139;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 140;
address_inb = 141;
data_ina = 16'hfffe;
data_inb = 16'h1;
#10;
address_ina = 142;
address_inb = 143;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 144;
address_inb = 145;
data_ina = 16'hfffe;
data_inb = 16'hfffe;
#10;
address_ina = 146;
address_inb = 147;
data_ina = 16'hffff;
data_inb = 16'h2;
#10;
address_ina = 148;
address_inb = 149;
data_ina = 16'hfffe;
data_inb = 16'h0;
#10;
address_ina = 150;
address_inb = 151;
data_ina = 16'h0;
data_inb = 16'hfffe;
#10;
address_ina = 152;
address_inb = 153;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 154;
address_inb = 155;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 156;
address_inb = 157;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 158;
address_inb = 159;
data_ina = 16'hfffe;
data_inb = 16'h0;
#10;
address_ina = 160;
address_inb = 161;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 162;
address_inb = 163;
data_ina = 16'h2;
data_inb = 16'h1;
#10;
address_ina = 164;
address_inb = 165;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 166;
address_inb = 167;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 168;
address_inb = 169;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 170;
address_inb = 171;
data_ina = 16'h0;
data_inb = 16'h2;
#10;
address_ina = 172;
address_inb = 173;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 174;
address_inb = 175;
data_ina = 16'h1;
data_inb = 16'h2;
#10;
address_ina = 176;
address_inb = 177;
data_ina = 16'h1;
data_inb = 16'h2;
#10;
address_ina = 178;
address_inb = 179;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 180;
address_inb = 181;
data_ina = 16'h0;
data_inb = 16'h3;
#10;
address_ina = 182;
address_inb = 183;
data_ina = 16'h3;
data_inb = 16'hffff;
#10;
address_ina = 184;
address_inb = 185;
data_ina = 16'h1;
data_inb = 16'h2;
#10;
address_ina = 186;
address_inb = 187;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 188;
address_inb = 189;
data_ina = 16'hfffe;
data_inb = 16'hfffe;
#10;
address_ina = 190;
address_inb = 191;
data_ina = 16'h1;
data_inb = 16'hfffe;
#10;
address_ina = 192;
address_inb = 193;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 194;
address_inb = 195;
data_ina = 16'h2;
data_inb = 16'h1;
#10;
address_ina = 196;
address_inb = 197;
data_ina = 16'hfffe;
data_inb = 16'hffff;
#10;
address_ina = 198;
address_inb = 199;
data_ina = 16'hfffe;
data_inb = 16'hfffd;
#10;
address_ina = 200;
address_inb = 201;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 202;
address_inb = 203;
data_ina = 16'h1;
data_inb = 16'hfffe;
#10;
address_ina = 204;
address_inb = 205;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 206;
address_inb = 207;
data_ina = 16'hffff;
data_inb = 16'hfffe;
#10;
address_ina = 208;
address_inb = 209;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 210;
address_inb = 211;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 212;
address_inb = 213;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 214;
address_inb = 215;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 216;
address_inb = 217;
data_ina = 16'h1;
data_inb = 16'hfffe;
#10;
address_ina = 218;
address_inb = 219;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 220;
address_inb = 221;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 222;
address_inb = 223;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 224;
address_inb = 225;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 226;
address_inb = 227;
data_ina = 16'hfffe;
data_inb = 16'h0;
#10;
address_ina = 228;
address_inb = 229;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 230;
address_inb = 231;
data_ina = 16'h0;
data_inb = 16'h2;
#10;
address_ina = 232;
address_inb = 233;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 234;
address_inb = 235;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 236;
address_inb = 237;
data_ina = 16'hffff;
data_inb = 16'hfffe;
#10;
address_ina = 238;
address_inb = 239;
data_ina = 16'h2;
data_inb = 16'h0;
#10;
address_ina = 240;
address_inb = 241;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 242;
address_inb = 243;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 244;
address_inb = 245;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 246;
address_inb = 247;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 248;
address_inb = 249;
data_ina = 16'h1;
data_inb = 16'h2;
#10;
address_ina = 250;
address_inb = 251;
data_ina = 16'h0;
data_inb = 16'hfffe;
#10;
address_ina = 252;
address_inb = 253;
data_ina = 16'hfffd;
data_inb = 16'h1;
#10;
address_ina = 254;
address_inb = 255;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
        wait(init_done);
        #30
        we = 0;
        // Start processing
         
		  #38000

        start = 0;



//        wait (wr_req);
//		  wait (!wr_req);
//		   rd_req = 1;
		  wait(done);
		  #20000
rd_req = 1;
        #70 
		  start = 1;
		 #80 
wait(rd_empty)
rd_req = 0;

$display("Finished the NTT test Number %d",test_num);
////Begin test number #22//////////////
rst = 1;

//#1000
start = 1;
mode = 0; //NTT 0 // INTT 1

// Reset for a few clock cycles

#1000

rst = 0;
test_num = test_num + 1;
#1000
we = 1;
address_ina = 0;
address_inb = 1;
data_ina = 16'hfffd;
data_inb = 16'h0;
#10;
address_ina = 2;
address_inb = 3;
data_ina = 16'h0;
data_inb = 16'h2;
#10;
address_ina = 4;
address_inb = 5;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 6;
address_inb = 7;
data_ina = 16'hffff;
data_inb = 16'h2;
#10;
address_ina = 8;
address_inb = 9;
data_ina = 16'h0;
data_inb = 16'hfffe;
#10;
address_ina = 10;
address_inb = 11;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 12;
address_inb = 13;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 14;
address_inb = 15;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 16;
address_inb = 17;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 18;
address_inb = 19;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 20;
address_inb = 21;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 22;
address_inb = 23;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 24;
address_inb = 25;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 26;
address_inb = 27;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 28;
address_inb = 29;
data_ina = 16'h2;
data_inb = 16'h0;
#10;
address_ina = 30;
address_inb = 31;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 32;
address_inb = 33;
data_ina = 16'h0;
data_inb = 16'h2;
#10;
address_ina = 34;
address_inb = 35;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 36;
address_inb = 37;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 38;
address_inb = 39;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 40;
address_inb = 41;
data_ina = 16'h0;
data_inb = 16'hfffe;
#10;
address_ina = 42;
address_inb = 43;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 44;
address_inb = 45;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 46;
address_inb = 47;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 48;
address_inb = 49;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 50;
address_inb = 51;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 52;
address_inb = 53;
data_ina = 16'h1;
data_inb = 16'hfffe;
#10;
address_ina = 54;
address_inb = 55;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 56;
address_inb = 57;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 58;
address_inb = 59;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 60;
address_inb = 61;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 62;
address_inb = 63;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 64;
address_inb = 65;
data_ina = 16'h1;
data_inb = 16'h2;
#10;
address_ina = 66;
address_inb = 67;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 68;
address_inb = 69;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 70;
address_inb = 71;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 72;
address_inb = 73;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 74;
address_inb = 75;
data_ina = 16'hfffe;
data_inb = 16'h1;
#10;
address_ina = 76;
address_inb = 77;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 78;
address_inb = 79;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 80;
address_inb = 81;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 82;
address_inb = 83;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 84;
address_inb = 85;
data_ina = 16'h2;
data_inb = 16'h2;
#10;
address_ina = 86;
address_inb = 87;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 88;
address_inb = 89;
data_ina = 16'h2;
data_inb = 16'hffff;
#10;
address_ina = 90;
address_inb = 91;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 92;
address_inb = 93;
data_ina = 16'h0;
data_inb = 16'h3;
#10;
address_ina = 94;
address_inb = 95;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 96;
address_inb = 97;
data_ina = 16'h2;
data_inb = 16'h0;
#10;
address_ina = 98;
address_inb = 99;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 100;
address_inb = 101;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 102;
address_inb = 103;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 104;
address_inb = 105;
data_ina = 16'hfffe;
data_inb = 16'h1;
#10;
address_ina = 106;
address_inb = 107;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 108;
address_inb = 109;
data_ina = 16'hfffe;
data_inb = 16'hfffe;
#10;
address_ina = 110;
address_inb = 111;
data_ina = 16'h1;
data_inb = 16'h2;
#10;
address_ina = 112;
address_inb = 113;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 114;
address_inb = 115;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 116;
address_inb = 117;
data_ina = 16'h2;
data_inb = 16'h0;
#10;
address_ina = 118;
address_inb = 119;
data_ina = 16'hfffe;
data_inb = 16'h1;
#10;
address_ina = 120;
address_inb = 121;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 122;
address_inb = 123;
data_ina = 16'hfffe;
data_inb = 16'hffff;
#10;
address_ina = 124;
address_inb = 125;
data_ina = 16'h3;
data_inb = 16'h1;
#10;
address_ina = 126;
address_inb = 127;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 128;
address_inb = 129;
data_ina = 16'hfffd;
data_inb = 16'h0;
#10;
address_ina = 130;
address_inb = 131;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 132;
address_inb = 133;
data_ina = 16'h0;
data_inb = 16'hfffe;
#10;
address_ina = 134;
address_inb = 135;
data_ina = 16'h1;
data_inb = 16'h2;
#10;
address_ina = 136;
address_inb = 137;
data_ina = 16'h2;
data_inb = 16'hffff;
#10;
address_ina = 138;
address_inb = 139;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 140;
address_inb = 141;
data_ina = 16'hfffe;
data_inb = 16'hffff;
#10;
address_ina = 142;
address_inb = 143;
data_ina = 16'h2;
data_inb = 16'h1;
#10;
address_ina = 144;
address_inb = 145;
data_ina = 16'h2;
data_inb = 16'h1;
#10;
address_ina = 146;
address_inb = 147;
data_ina = 16'hfffe;
data_inb = 16'h0;
#10;
address_ina = 148;
address_inb = 149;
data_ina = 16'h1;
data_inb = 16'h2;
#10;
address_ina = 150;
address_inb = 151;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 152;
address_inb = 153;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 154;
address_inb = 155;
data_ina = 16'h2;
data_inb = 16'hffff;
#10;
address_ina = 156;
address_inb = 157;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 158;
address_inb = 159;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 160;
address_inb = 161;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 162;
address_inb = 163;
data_ina = 16'h2;
data_inb = 16'h0;
#10;
address_ina = 164;
address_inb = 165;
data_ina = 16'hffff;
data_inb = 16'h2;
#10;
address_ina = 166;
address_inb = 167;
data_ina = 16'h0;
data_inb = 16'h2;
#10;
address_ina = 168;
address_inb = 169;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 170;
address_inb = 171;
data_ina = 16'h3;
data_inb = 16'h0;
#10;
address_ina = 172;
address_inb = 173;
data_ina = 16'h1;
data_inb = 16'h2;
#10;
address_ina = 174;
address_inb = 175;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 176;
address_inb = 177;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 178;
address_inb = 179;
data_ina = 16'hfffe;
data_inb = 16'h2;
#10;
address_ina = 180;
address_inb = 181;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 182;
address_inb = 183;
data_ina = 16'h1;
data_inb = 16'h2;
#10;
address_ina = 184;
address_inb = 185;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 186;
address_inb = 187;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 188;
address_inb = 189;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 190;
address_inb = 191;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 192;
address_inb = 193;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 194;
address_inb = 195;
data_ina = 16'hfffe;
data_inb = 16'h0;
#10;
address_ina = 196;
address_inb = 197;
data_ina = 16'hfffe;
data_inb = 16'h1;
#10;
address_ina = 198;
address_inb = 199;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 200;
address_inb = 201;
data_ina = 16'hfffe;
data_inb = 16'h0;
#10;
address_ina = 202;
address_inb = 203;
data_ina = 16'hfffd;
data_inb = 16'h0;
#10;
address_ina = 204;
address_inb = 205;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 206;
address_inb = 207;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 208;
address_inb = 209;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 210;
address_inb = 211;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 212;
address_inb = 213;
data_ina = 16'h0;
data_inb = 16'h2;
#10;
address_ina = 214;
address_inb = 215;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 216;
address_inb = 217;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 218;
address_inb = 219;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 220;
address_inb = 221;
data_ina = 16'hffff;
data_inb = 16'hfffe;
#10;
address_ina = 222;
address_inb = 223;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 224;
address_inb = 225;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 226;
address_inb = 227;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 228;
address_inb = 229;
data_ina = 16'hfffe;
data_inb = 16'h1;
#10;
address_ina = 230;
address_inb = 231;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 232;
address_inb = 233;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 234;
address_inb = 235;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 236;
address_inb = 237;
data_ina = 16'hffff;
data_inb = 16'hfffe;
#10;
address_ina = 238;
address_inb = 239;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 240;
address_inb = 241;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 242;
address_inb = 243;
data_ina = 16'h2;
data_inb = 16'hfffe;
#10;
address_ina = 244;
address_inb = 245;
data_ina = 16'hfffe;
data_inb = 16'hffff;
#10;
address_ina = 246;
address_inb = 247;
data_ina = 16'h2;
data_inb = 16'h2;
#10;
address_ina = 248;
address_inb = 249;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 250;
address_inb = 251;
data_ina = 16'hfffe;
data_inb = 16'h0;
#10;
address_ina = 252;
address_inb = 253;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 254;
address_inb = 255;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
        wait(init_done);
        #30
        we = 0;
        // Start processing
         
		  #38000

        start = 0;



//        wait (wr_req);
//		  wait (!wr_req);
//		   rd_req = 1;
		  wait(done);
		  #20000
rd_req = 1;
        #70 
		  start = 1;
		 #80 
wait(rd_empty)
rd_req = 0;

$display("Finished the NTT test Number %d",test_num);
////Begin test number #23//////////////
rst = 1;

//#1000
start = 1;
mode = 1; //NTT 0 // INTT 1

// Reset for a few clock cycles

#1000

rst = 0;
test_num = test_num + 1;
#1000
we = 1;
address_ina = 0;
address_inb = 1;
data_ina = 16'he2;
data_inb = 16'h583;
#10;
address_ina = 2;
address_inb = 3;
data_ina = 16'hfc89;
data_inb = 16'h7d;
#10;
address_ina = 4;
address_inb = 5;
data_ina = 16'hfdfe;
data_inb = 16'h25e;
#10;
address_ina = 6;
address_inb = 7;
data_ina = 16'h677;
data_inb = 16'hfb65;
#10;
address_ina = 8;
address_inb = 9;
data_ina = 16'h29d;
data_inb = 16'hff07;
#10;
address_ina = 10;
address_inb = 11;
data_ina = 16'h64e;
data_inb = 16'hff6e;
#10;
address_ina = 12;
address_inb = 13;
data_ina = 16'h7e;
data_inb = 16'hff2b;
#10;
address_ina = 14;
address_inb = 15;
data_ina = 16'hfd32;
data_inb = 16'h420;
#10;
address_ina = 16;
address_inb = 17;
data_ina = 16'hf985;
data_inb = 16'h26f;
#10;
address_ina = 18;
address_inb = 19;
data_ina = 16'hfd48;
data_inb = 16'hfa4b;
#10;
address_ina = 20;
address_inb = 21;
data_ina = 16'h5c0;
data_inb = 16'h299;
#10;
address_ina = 22;
address_inb = 23;
data_ina = 16'h2c1;
data_inb = 16'hfda1;
#10;
address_ina = 24;
address_inb = 25;
data_ina = 16'h33b;
data_inb = 16'h628;
#10;
address_ina = 26;
address_inb = 27;
data_ina = 16'hfe0e;
data_inb = 16'hf9fc;
#10;
address_ina = 28;
address_inb = 29;
data_ina = 16'hfd1e;
data_inb = 16'h11;
#10;
address_ina = 30;
address_inb = 31;
data_ina = 16'h554;
data_inb = 16'hfbc6;
#10;
address_ina = 32;
address_inb = 33;
data_ina = 16'h36a;
data_inb = 16'hfa62;
#10;
address_ina = 34;
address_inb = 35;
data_ina = 16'hf98c;
data_inb = 16'h269;
#10;
address_ina = 36;
address_inb = 37;
data_ina = 16'hfb14;
data_inb = 16'h40a;
#10;
address_ina = 38;
address_inb = 39;
data_ina = 16'h5e8;
data_inb = 16'h2fa;
#10;
address_ina = 40;
address_inb = 41;
data_ina = 16'hdb;
data_inb = 16'hfc80;
#10;
address_ina = 42;
address_inb = 43;
data_ina = 16'h26f;
data_inb = 16'h470;
#10;
address_ina = 44;
address_inb = 45;
data_ina = 16'h3;
data_inb = 16'hfd06;
#10;
address_ina = 46;
address_inb = 47;
data_ina = 16'h467;
data_inb = 16'hfe7e;
#10;
address_ina = 48;
address_inb = 49;
data_ina = 16'hfef2;
data_inb = 16'hff7d;
#10;
address_ina = 50;
address_inb = 51;
data_ina = 16'hff56;
data_inb = 16'hfd4b;
#10;
address_ina = 52;
address_inb = 53;
data_ina = 16'h272;
data_inb = 16'hffba;
#10;
address_ina = 54;
address_inb = 55;
data_ina = 16'hfd9b;
data_inb = 16'hfeef;
#10;
address_ina = 56;
address_inb = 57;
data_ina = 16'hfce8;
data_inb = 16'hfc9a;
#10;
address_ina = 58;
address_inb = 59;
data_ina = 16'h45e;
data_inb = 16'hfc4d;
#10;
address_ina = 60;
address_inb = 61;
data_ina = 16'h55a;
data_inb = 16'hfd10;
#10;
address_ina = 62;
address_inb = 63;
data_ina = 16'hfdef;
data_inb = 16'hfb13;
#10;
address_ina = 64;
address_inb = 65;
data_ina = 16'h528;
data_inb = 16'h1a1;
#10;
address_ina = 66;
address_inb = 67;
data_ina = 16'hfb8f;
data_inb = 16'h114;
#10;
address_ina = 68;
address_inb = 69;
data_ina = 16'h4b5;
data_inb = 16'h192;
#10;
address_ina = 70;
address_inb = 71;
data_ina = 16'hff2a;
data_inb = 16'hffe7;
#10;
address_ina = 72;
address_inb = 73;
data_ina = 16'hf994;
data_inb = 16'h104;
#10;
address_ina = 74;
address_inb = 75;
data_ina = 16'hf9e0;
data_inb = 16'h557;
#10;
address_ina = 76;
address_inb = 77;
data_ina = 16'h4c7;
data_inb = 16'h288;
#10;
address_ina = 78;
address_inb = 79;
data_ina = 16'hfadd;
data_inb = 16'h55;
#10;
address_ina = 80;
address_inb = 81;
data_ina = 16'hf9d9;
data_inb = 16'hfa71;
#10;
address_ina = 82;
address_inb = 83;
data_ina = 16'h4fa;
data_inb = 16'h0;
#10;
address_ina = 84;
address_inb = 85;
data_ina = 16'ha5;
data_inb = 16'hfcb7;
#10;
address_ina = 86;
address_inb = 87;
data_ina = 16'h178;
data_inb = 16'hfe3b;
#10;
address_ina = 88;
address_inb = 89;
data_ina = 16'h57b;
data_inb = 16'h4dd;
#10;
address_ina = 90;
address_inb = 91;
data_ina = 16'h58c;
data_inb = 16'hfe95;
#10;
address_ina = 92;
address_inb = 93;
data_ina = 16'hfc94;
data_inb = 16'h37;
#10;
address_ina = 94;
address_inb = 95;
data_ina = 16'hfa42;
data_inb = 16'hfb93;
#10;
address_ina = 96;
address_inb = 97;
data_ina = 16'hff02;
data_inb = 16'h243;
#10;
address_ina = 98;
address_inb = 99;
data_ina = 16'h3d5;
data_inb = 16'h43f;
#10;
address_ina = 100;
address_inb = 101;
data_ina = 16'h3fc;
data_inb = 16'hf9de;
#10;
address_ina = 102;
address_inb = 103;
data_ina = 16'h483;
data_inb = 16'h55;
#10;
address_ina = 104;
address_inb = 105;
data_ina = 16'h3c9;
data_inb = 16'hf9c3;
#10;
address_ina = 106;
address_inb = 107;
data_ina = 16'h56c;
data_inb = 16'h45c;
#10;
address_ina = 108;
address_inb = 109;
data_ina = 16'hfecb;
data_inb = 16'h542;
#10;
address_ina = 110;
address_inb = 111;
data_ina = 16'hfed8;
data_inb = 16'hfad8;
#10;
address_ina = 112;
address_inb = 113;
data_ina = 16'hfb79;
data_inb = 16'h3a;
#10;
address_ina = 114;
address_inb = 115;
data_ina = 16'hfec4;
data_inb = 16'hff31;
#10;
address_ina = 116;
address_inb = 117;
data_ina = 16'h153;
data_inb = 16'h491;
#10;
address_ina = 118;
address_inb = 119;
data_ina = 16'h49f;
data_inb = 16'h50e;
#10;
address_ina = 120;
address_inb = 121;
data_ina = 16'he8;
data_inb = 16'h524;
#10;
address_ina = 122;
address_inb = 123;
data_ina = 16'hfdc8;
data_inb = 16'hf9c3;
#10;
address_ina = 124;
address_inb = 125;
data_ina = 16'hffa8;
data_inb = 16'h23d;
#10;
address_ina = 126;
address_inb = 127;
data_ina = 16'h316;
data_inb = 16'hfdbb;
#10;
address_ina = 128;
address_inb = 129;
data_ina = 16'hfeb3;
data_inb = 16'hfcfa;
#10;
address_ina = 130;
address_inb = 131;
data_ina = 16'h22;
data_inb = 16'hfaf4;
#10;
address_ina = 132;
address_inb = 133;
data_ina = 16'hff3c;
data_inb = 16'hfa0b;
#10;
address_ina = 134;
address_inb = 135;
data_ina = 16'hfcde;
data_inb = 16'h27e;
#10;
address_ina = 136;
address_inb = 137;
data_ina = 16'hfd18;
data_inb = 16'h286;
#10;
address_ina = 138;
address_inb = 139;
data_ina = 16'hfc1d;
data_inb = 16'h4f0;
#10;
address_ina = 140;
address_inb = 141;
data_ina = 16'h399;
data_inb = 16'hfa35;
#10;
address_ina = 142;
address_inb = 143;
data_ina = 16'hfc9e;
data_inb = 16'hf98f;
#10;
address_ina = 144;
address_inb = 145;
data_ina = 16'hfdd2;
data_inb = 16'hfbf9;
#10;
address_ina = 146;
address_inb = 147;
data_ina = 16'h110;
data_inb = 16'h349;
#10;
address_ina = 148;
address_inb = 149;
data_ina = 16'hfc14;
data_inb = 16'h4fb;
#10;
address_ina = 150;
address_inb = 151;
data_ina = 16'h5af;
data_inb = 16'hffb3;
#10;
address_ina = 152;
address_inb = 153;
data_ina = 16'hfc4f;
data_inb = 16'hf983;
#10;
address_ina = 154;
address_inb = 155;
data_ina = 16'hfa18;
data_inb = 16'hfde4;
#10;
address_ina = 156;
address_inb = 157;
data_ina = 16'hf2;
data_inb = 16'hfa43;
#10;
address_ina = 158;
address_inb = 159;
data_ina = 16'h5a1;
data_inb = 16'hfa76;
#10;
address_ina = 160;
address_inb = 161;
data_ina = 16'h5ac;
data_inb = 16'hff33;
#10;
address_ina = 162;
address_inb = 163;
data_ina = 16'hfacb;
data_inb = 16'hfbe6;
#10;
address_ina = 164;
address_inb = 165;
data_ina = 16'hfaf3;
data_inb = 16'hfa69;
#10;
address_ina = 166;
address_inb = 167;
data_ina = 16'hfe81;
data_inb = 16'h51d;
#10;
address_ina = 168;
address_inb = 169;
data_ina = 16'h12d;
data_inb = 16'h46e;
#10;
address_ina = 170;
address_inb = 171;
data_ina = 16'hfa20;
data_inb = 16'hfc44;
#10;
address_ina = 172;
address_inb = 173;
data_ina = 16'h3e6;
data_inb = 16'hfae6;
#10;
address_ina = 174;
address_inb = 175;
data_ina = 16'h107;
data_inb = 16'h143;
#10;
address_ina = 176;
address_inb = 177;
data_ina = 16'hfa11;
data_inb = 16'hfb4d;
#10;
address_ina = 178;
address_inb = 179;
data_ina = 16'hac;
data_inb = 16'h66f;
#10;
address_ina = 180;
address_inb = 181;
data_ina = 16'h124;
data_inb = 16'h285;
#10;
address_ina = 182;
address_inb = 183;
data_ina = 16'hff02;
data_inb = 16'h4f4;
#10;
address_ina = 184;
address_inb = 185;
data_ina = 16'hfc78;
data_inb = 16'hfb4a;
#10;
address_ina = 186;
address_inb = 187;
data_ina = 16'hff6d;
data_inb = 16'h1b2;
#10;
address_ina = 188;
address_inb = 189;
data_ina = 16'h3de;
data_inb = 16'h47d;
#10;
address_ina = 190;
address_inb = 191;
data_ina = 16'h362;
data_inb = 16'h5f6;
#10;
address_ina = 192;
address_inb = 193;
data_ina = 16'hfd13;
data_inb = 16'hfd91;
#10;
address_ina = 194;
address_inb = 195;
data_ina = 16'h302;
data_inb = 16'h1bd;
#10;
address_ina = 196;
address_inb = 197;
data_ina = 16'h2a0;
data_inb = 16'hf9ec;
#10;
address_ina = 198;
address_inb = 199;
data_ina = 16'h2fd;
data_inb = 16'hfaec;
#10;
address_ina = 200;
address_inb = 201;
data_ina = 16'hf98d;
data_inb = 16'hf9a0;
#10;
address_ina = 202;
address_inb = 203;
data_ina = 16'hf996;
data_inb = 16'hfb7f;
#10;
address_ina = 204;
address_inb = 205;
data_ina = 16'hfbcf;
data_inb = 16'h3b3;
#10;
address_ina = 206;
address_inb = 207;
data_ina = 16'hff78;
data_inb = 16'h5d1;
#10;
address_ina = 208;
address_inb = 209;
data_ina = 16'h2e;
data_inb = 16'hfdc8;
#10;
address_ina = 210;
address_inb = 211;
data_ina = 16'hfda2;
data_inb = 16'h3fa;
#10;
address_ina = 212;
address_inb = 213;
data_ina = 16'hf9b2;
data_inb = 16'hfdc6;
#10;
address_ina = 214;
address_inb = 215;
data_ina = 16'h2d2;
data_inb = 16'h4cb;
#10;
address_ina = 216;
address_inb = 217;
data_ina = 16'hf9d2;
data_inb = 16'h2ed;
#10;
address_ina = 218;
address_inb = 219;
data_ina = 16'hfeb2;
data_inb = 16'hfdf8;
#10;
address_ina = 220;
address_inb = 221;
data_ina = 16'hff24;
data_inb = 16'hfbd5;
#10;
address_ina = 222;
address_inb = 223;
data_ina = 16'hfa61;
data_inb = 16'h1eb;
#10;
address_ina = 224;
address_inb = 225;
data_ina = 16'hff14;
data_inb = 16'h49b;
#10;
address_ina = 226;
address_inb = 227;
data_ina = 16'hfd8c;
data_inb = 16'hf9fa;
#10;
address_ina = 228;
address_inb = 229;
data_ina = 16'hfeb6;
data_inb = 16'hfb29;
#10;
address_ina = 230;
address_inb = 231;
data_ina = 16'hff46;
data_inb = 16'h59f;
#10;
address_ina = 232;
address_inb = 233;
data_ina = 16'h443;
data_inb = 16'h21a;
#10;
address_ina = 234;
address_inb = 235;
data_ina = 16'hff97;
data_inb = 16'h365;
#10;
address_ina = 236;
address_inb = 237;
data_ina = 16'hfbec;
data_inb = 16'h235;
#10;
address_ina = 238;
address_inb = 239;
data_ina = 16'h529;
data_inb = 16'h48b;
#10;
address_ina = 240;
address_inb = 241;
data_ina = 16'h22f;
data_inb = 16'hf9c4;
#10;
address_ina = 242;
address_inb = 243;
data_ina = 16'h37;
data_inb = 16'hfccb;
#10;
address_ina = 244;
address_inb = 245;
data_ina = 16'hfcf4;
data_inb = 16'hfb08;
#10;
address_ina = 246;
address_inb = 247;
data_ina = 16'h1f1;
data_inb = 16'h544;
#10;
address_ina = 248;
address_inb = 249;
data_ina = 16'hfd28;
data_inb = 16'h653;
#10;
address_ina = 250;
address_inb = 251;
data_ina = 16'hff03;
data_inb = 16'hfd9b;
#10;
address_ina = 252;
address_inb = 253;
data_ina = 16'hfc77;
data_inb = 16'h202;
#10;
address_ina = 254;
address_inb = 255;
data_ina = 16'hfa80;
data_inb = 16'h1e8;
#10;
        wait(init_done);
        #30
        we = 0;
        // Start processing
         
		  #38000

        start = 0;



//        wait (wr_req);
//		  wait (!wr_req);
//		   rd_req = 1;
		  wait(done);
		  #20000
rd_req = 1;
        #70 
		  start = 1;
		 #80 
wait(rd_empty)
rd_req = 0;

$display("Finished the NTT test Number %d",test_num);
////Begin test number #24//////////////
rst = 1;

//#1000
start = 1;
mode = 1; //NTT 0 // INTT 1

// Reset for a few clock cycles

#1000

rst = 0;
test_num = test_num + 1;
#1000
we = 1;
address_ina = 0;
address_inb = 1;
data_ina = 16'h128;
data_inb = 16'hff6e;
#10;
address_ina = 2;
address_inb = 3;
data_ina = 16'hfad8;
data_inb = 16'h3c8;
#10;
address_ina = 4;
address_inb = 5;
data_ina = 16'h475;
data_inb = 16'hff88;
#10;
address_ina = 6;
address_inb = 7;
data_ina = 16'h3c4;
data_inb = 16'h3de;
#10;
address_ina = 8;
address_inb = 9;
data_ina = 16'hff64;
data_inb = 16'hf992;
#10;
address_ina = 10;
address_inb = 11;
data_ina = 16'hfd45;
data_inb = 16'h607;
#10;
address_ina = 12;
address_inb = 13;
data_ina = 16'h5b9;
data_inb = 16'hfa5e;
#10;
address_ina = 14;
address_inb = 15;
data_ina = 16'h424;
data_inb = 16'h473;
#10;
address_ina = 16;
address_inb = 17;
data_ina = 16'hfdc3;
data_inb = 16'hfe59;
#10;
address_ina = 18;
address_inb = 19;
data_ina = 16'h308;
data_inb = 16'hfccc;
#10;
address_ina = 20;
address_inb = 21;
data_ina = 16'hfad2;
data_inb = 16'hfe85;
#10;
address_ina = 22;
address_inb = 23;
data_ina = 16'hfbc0;
data_inb = 16'hffc6;
#10;
address_ina = 24;
address_inb = 25;
data_ina = 16'hfb91;
data_inb = 16'hfc05;
#10;
address_ina = 26;
address_inb = 27;
data_ina = 16'hf9a2;
data_inb = 16'h2b5;
#10;
address_ina = 28;
address_inb = 29;
data_ina = 16'hfb34;
data_inb = 16'h5ca;
#10;
address_ina = 30;
address_inb = 31;
data_ina = 16'hfe87;
data_inb = 16'h40e;
#10;
address_ina = 32;
address_inb = 33;
data_ina = 16'hfc2f;
data_inb = 16'h50c;
#10;
address_ina = 34;
address_inb = 35;
data_ina = 16'hfcdb;
data_inb = 16'h1c2;
#10;
address_ina = 36;
address_inb = 37;
data_ina = 16'hff5e;
data_inb = 16'hf9bc;
#10;
address_ina = 38;
address_inb = 39;
data_ina = 16'hfca9;
data_inb = 16'h2b;
#10;
address_ina = 40;
address_inb = 41;
data_ina = 16'hfdf3;
data_inb = 16'h629;
#10;
address_ina = 42;
address_inb = 43;
data_ina = 16'h566;
data_inb = 16'hfe74;
#10;
address_ina = 44;
address_inb = 45;
data_ina = 16'hfed4;
data_inb = 16'h28c;
#10;
address_ina = 46;
address_inb = 47;
data_ina = 16'hfea6;
data_inb = 16'hfaed;
#10;
address_ina = 48;
address_inb = 49;
data_ina = 16'h2f3;
data_inb = 16'hdc;
#10;
address_ina = 50;
address_inb = 51;
data_ina = 16'h5cd;
data_inb = 16'hfbba;
#10;
address_ina = 52;
address_inb = 53;
data_ina = 16'hfabc;
data_inb = 16'hfabf;
#10;
address_ina = 54;
address_inb = 55;
data_ina = 16'hca;
data_inb = 16'h3db;
#10;
address_ina = 56;
address_inb = 57;
data_ina = 16'h62b;
data_inb = 16'h55b;
#10;
address_ina = 58;
address_inb = 59;
data_ina = 16'h5c7;
data_inb = 16'h2f;
#10;
address_ina = 60;
address_inb = 61;
data_ina = 16'h1d2;
data_inb = 16'h2af;
#10;
address_ina = 62;
address_inb = 63;
data_ina = 16'hfdd9;
data_inb = 16'hfb35;
#10;
address_ina = 64;
address_inb = 65;
data_ina = 16'hfa2c;
data_inb = 16'h27a;
#10;
address_ina = 66;
address_inb = 67;
data_ina = 16'hfbb4;
data_inb = 16'h4a5;
#10;
address_ina = 68;
address_inb = 69;
data_ina = 16'hfb57;
data_inb = 16'hfc40;
#10;
address_ina = 70;
address_inb = 71;
data_ina = 16'hfffa;
data_inb = 16'hf98c;
#10;
address_ina = 72;
address_inb = 73;
data_ina = 16'h5b6;
data_inb = 16'h529;
#10;
address_ina = 74;
address_inb = 75;
data_ina = 16'h1d;
data_inb = 16'h274;
#10;
address_ina = 76;
address_inb = 77;
data_ina = 16'hff69;
data_inb = 16'h322;
#10;
address_ina = 78;
address_inb = 79;
data_ina = 16'hfb01;
data_inb = 16'hff7f;
#10;
address_ina = 80;
address_inb = 81;
data_ina = 16'hf9a1;
data_inb = 16'hfea0;
#10;
address_ina = 82;
address_inb = 83;
data_ina = 16'hfac3;
data_inb = 16'h2ce;
#10;
address_ina = 84;
address_inb = 85;
data_ina = 16'h658;
data_inb = 16'hfbeb;
#10;
address_ina = 86;
address_inb = 87;
data_ina = 16'h58e;
data_inb = 16'h23a;
#10;
address_ina = 88;
address_inb = 89;
data_ina = 16'h93;
data_inb = 16'h24;
#10;
address_ina = 90;
address_inb = 91;
data_ina = 16'h42d;
data_inb = 16'hfcbf;
#10;
address_ina = 92;
address_inb = 93;
data_ina = 16'hfb74;
data_inb = 16'hfea0;
#10;
address_ina = 94;
address_inb = 95;
data_ina = 16'hfe9e;
data_inb = 16'hfb7e;
#10;
address_ina = 96;
address_inb = 97;
data_ina = 16'hffa9;
data_inb = 16'h3a7;
#10;
address_ina = 98;
address_inb = 99;
data_ina = 16'hf98d;
data_inb = 16'hfecb;
#10;
address_ina = 100;
address_inb = 101;
data_ina = 16'hfcd8;
data_inb = 16'hfdff;
#10;
address_ina = 102;
address_inb = 103;
data_ina = 16'hfff5;
data_inb = 16'hffce;
#10;
address_ina = 104;
address_inb = 105;
data_ina = 16'hfa8e;
data_inb = 16'hfe28;
#10;
address_ina = 106;
address_inb = 107;
data_ina = 16'h5ef;
data_inb = 16'hfc26;
#10;
address_ina = 108;
address_inb = 109;
data_ina = 16'h349;
data_inb = 16'hf9f9;
#10;
address_ina = 110;
address_inb = 111;
data_ina = 16'hfd78;
data_inb = 16'hfdfc;
#10;
address_ina = 112;
address_inb = 113;
data_ina = 16'hfe74;
data_inb = 16'h66f;
#10;
address_ina = 114;
address_inb = 115;
data_ina = 16'h58c;
data_inb = 16'hfce9;
#10;
address_ina = 116;
address_inb = 117;
data_ina = 16'h339;
data_inb = 16'hfe74;
#10;
address_ina = 118;
address_inb = 119;
data_ina = 16'hfd2e;
data_inb = 16'hf98f;
#10;
address_ina = 120;
address_inb = 121;
data_ina = 16'hfb73;
data_inb = 16'hee;
#10;
address_ina = 122;
address_inb = 123;
data_ina = 16'h13e;
data_inb = 16'hfbef;
#10;
address_ina = 124;
address_inb = 125;
data_ina = 16'h3c7;
data_inb = 16'hfec7;
#10;
address_ina = 126;
address_inb = 127;
data_ina = 16'h253;
data_inb = 16'hfbac;
#10;
address_ina = 128;
address_inb = 129;
data_ina = 16'hffdc;
data_inb = 16'hfc1c;
#10;
address_ina = 130;
address_inb = 131;
data_ina = 16'hfefa;
data_inb = 16'h21d;
#10;
address_ina = 132;
address_inb = 133;
data_ina = 16'h5e1;
data_inb = 16'hfa95;
#10;
address_ina = 134;
address_inb = 135;
data_ina = 16'h24a;
data_inb = 16'hfbb1;
#10;
address_ina = 136;
address_inb = 137;
data_ina = 16'h63e;
data_inb = 16'hff5b;
#10;
address_ina = 138;
address_inb = 139;
data_ina = 16'hfd3b;
data_inb = 16'hfe69;
#10;
address_ina = 140;
address_inb = 141;
data_ina = 16'h49f;
data_inb = 16'hf98a;
#10;
address_ina = 142;
address_inb = 143;
data_ina = 16'hfd0c;
data_inb = 16'hfcf2;
#10;
address_ina = 144;
address_inb = 145;
data_ina = 16'h5ef;
data_inb = 16'hfee5;
#10;
address_ina = 146;
address_inb = 147;
data_ina = 16'h4c1;
data_inb = 16'h219;
#10;
address_ina = 148;
address_inb = 149;
data_ina = 16'h81;
data_inb = 16'h36c;
#10;
address_ina = 150;
address_inb = 151;
data_ina = 16'h19a;
data_inb = 16'h38f;
#10;
address_ina = 152;
address_inb = 153;
data_ina = 16'hfd6d;
data_inb = 16'hfa1d;
#10;
address_ina = 154;
address_inb = 155;
data_ina = 16'h44c;
data_inb = 16'h5fa;
#10;
address_ina = 156;
address_inb = 157;
data_ina = 16'hfa12;
data_inb = 16'h512;
#10;
address_ina = 158;
address_inb = 159;
data_ina = 16'h31a;
data_inb = 16'hfb0f;
#10;
address_ina = 160;
address_inb = 161;
data_ina = 16'h1d0;
data_inb = 16'hfe48;
#10;
address_ina = 162;
address_inb = 163;
data_ina = 16'h1c7;
data_inb = 16'hfc55;
#10;
address_ina = 164;
address_inb = 165;
data_ina = 16'h4de;
data_inb = 16'hc2;
#10;
address_ina = 166;
address_inb = 167;
data_ina = 16'hfa10;
data_inb = 16'hfff5;
#10;
address_ina = 168;
address_inb = 169;
data_ina = 16'hff75;
data_inb = 16'hffa4;
#10;
address_ina = 170;
address_inb = 171;
data_ina = 16'h46c;
data_inb = 16'hfdcc;
#10;
address_ina = 172;
address_inb = 173;
data_ina = 16'h532;
data_inb = 16'hff4e;
#10;
address_ina = 174;
address_inb = 175;
data_ina = 16'hfd44;
data_inb = 16'h33f;
#10;
address_ina = 176;
address_inb = 177;
data_ina = 16'h4d8;
data_inb = 16'hfd6c;
#10;
address_ina = 178;
address_inb = 179;
data_ina = 16'h1e5;
data_inb = 16'hfb36;
#10;
address_ina = 180;
address_inb = 181;
data_ina = 16'h5a1;
data_inb = 16'hfe3d;
#10;
address_ina = 182;
address_inb = 183;
data_ina = 16'hfce5;
data_inb = 16'h36;
#10;
address_ina = 184;
address_inb = 185;
data_ina = 16'h3ff;
data_inb = 16'hfcf7;
#10;
address_ina = 186;
address_inb = 187;
data_ina = 16'h494;
data_inb = 16'hfa8e;
#10;
address_ina = 188;
address_inb = 189;
data_ina = 16'h35d;
data_inb = 16'hffac;
#10;
address_ina = 190;
address_inb = 191;
data_ina = 16'hfec7;
data_inb = 16'h635;
#10;
address_ina = 192;
address_inb = 193;
data_ina = 16'h164;
data_inb = 16'h4c4;
#10;
address_ina = 194;
address_inb = 195;
data_ina = 16'h430;
data_inb = 16'hfa55;
#10;
address_ina = 196;
address_inb = 197;
data_ina = 16'hfc96;
data_inb = 16'hffd6;
#10;
address_ina = 198;
address_inb = 199;
data_ina = 16'hfebd;
data_inb = 16'h34;
#10;
address_ina = 200;
address_inb = 201;
data_ina = 16'hfd16;
data_inb = 16'h247;
#10;
address_ina = 202;
address_inb = 203;
data_ina = 16'hfa92;
data_inb = 16'hf99f;
#10;
address_ina = 204;
address_inb = 205;
data_ina = 16'h116;
data_inb = 16'hff8b;
#10;
address_ina = 206;
address_inb = 207;
data_ina = 16'hfc0f;
data_inb = 16'he6;
#10;
address_ina = 208;
address_inb = 209;
data_ina = 16'hfb4a;
data_inb = 16'h585;
#10;
address_ina = 210;
address_inb = 211;
data_ina = 16'h21;
data_inb = 16'h2f2;
#10;
address_ina = 212;
address_inb = 213;
data_ina = 16'hfc20;
data_inb = 16'hff2b;
#10;
address_ina = 214;
address_inb = 215;
data_ina = 16'h4dd;
data_inb = 16'hfc86;
#10;
address_ina = 216;
address_inb = 217;
data_ina = 16'h1f1;
data_inb = 16'h22;
#10;
address_ina = 218;
address_inb = 219;
data_ina = 16'hfbcf;
data_inb = 16'hfa03;
#10;
address_ina = 220;
address_inb = 221;
data_ina = 16'h5f;
data_inb = 16'hfb65;
#10;
address_ina = 222;
address_inb = 223;
data_ina = 16'h4d6;
data_inb = 16'h19c;
#10;
address_ina = 224;
address_inb = 225;
data_ina = 16'h15d;
data_inb = 16'h29c;
#10;
address_ina = 226;
address_inb = 227;
data_ina = 16'hf9ba;
data_inb = 16'hfbf9;
#10;
address_ina = 228;
address_inb = 229;
data_ina = 16'hfe88;
data_inb = 16'hffd8;
#10;
address_ina = 230;
address_inb = 231;
data_ina = 16'h78;
data_inb = 16'hfc6f;
#10;
address_ina = 232;
address_inb = 233;
data_ina = 16'h346;
data_inb = 16'hfe07;
#10;
address_ina = 234;
address_inb = 235;
data_ina = 16'hfdc7;
data_inb = 16'hffa9;
#10;
address_ina = 236;
address_inb = 237;
data_ina = 16'h2c5;
data_inb = 16'hff11;
#10;
address_ina = 238;
address_inb = 239;
data_ina = 16'h573;
data_inb = 16'h1e2;
#10;
address_ina = 240;
address_inb = 241;
data_ina = 16'hff6f;
data_inb = 16'h1ed;
#10;
address_ina = 242;
address_inb = 243;
data_ina = 16'hfe7a;
data_inb = 16'h45f;
#10;
address_ina = 244;
address_inb = 245;
data_ina = 16'hfc40;
data_inb = 16'h4df;
#10;
address_ina = 246;
address_inb = 247;
data_ina = 16'hfd0a;
data_inb = 16'hff4e;
#10;
address_ina = 248;
address_inb = 249;
data_ina = 16'hfca7;
data_inb = 16'h18;
#10;
address_ina = 250;
address_inb = 251;
data_ina = 16'hff7b;
data_inb = 16'he7;
#10;
address_ina = 252;
address_inb = 253;
data_ina = 16'hfc;
data_inb = 16'h613;
#10;
address_ina = 254;
address_inb = 255;
data_ina = 16'h4c5;
data_inb = 16'h57;
#10;
        wait(init_done);
        #30
        we = 0;
        // Start processing
         
		  #38000

        start = 0;



//        wait (wr_req);
//		  wait (!wr_req);
//		   rd_req = 1;
		  wait(done);
		  #20000
rd_req = 1;
        #70 
		  start = 1;
		 #80 
wait(rd_empty)
rd_req = 0;

$display("Finished the NTT test Number %d",test_num);
////Begin test number #25//////////////
rst = 1;

//#1000
start = 1;
mode = 1; //NTT 0 // INTT 1

// Reset for a few clock cycles

#1000

rst = 0;
test_num = test_num + 1;
#1000
we = 1;
address_ina = 0;
address_inb = 1;
data_ina = 16'hfc76;
data_inb = 16'h43;
#10;
address_ina = 2;
address_inb = 3;
data_ina = 16'hf98a;
data_inb = 16'h46a;
#10;
address_ina = 4;
address_inb = 5;
data_ina = 16'h283;
data_inb = 16'hfd;
#10;
address_ina = 6;
address_inb = 7;
data_ina = 16'hfbea;
data_inb = 16'hff4c;
#10;
address_ina = 8;
address_inb = 9;
data_ina = 16'hfce2;
data_inb = 16'hfe15;
#10;
address_ina = 10;
address_inb = 11;
data_ina = 16'hef;
data_inb = 16'h607;
#10;
address_ina = 12;
address_inb = 13;
data_ina = 16'hfc16;
data_inb = 16'hfbb6;
#10;
address_ina = 14;
address_inb = 15;
data_ina = 16'h4c6;
data_inb = 16'hfc9b;
#10;
address_ina = 16;
address_inb = 17;
data_ina = 16'h20b;
data_inb = 16'h128;
#10;
address_ina = 18;
address_inb = 19;
data_ina = 16'hffec;
data_inb = 16'h26c;
#10;
address_ina = 20;
address_inb = 21;
data_ina = 16'hff93;
data_inb = 16'hfc18;
#10;
address_ina = 22;
address_inb = 23;
data_ina = 16'h54a;
data_inb = 16'hfcc8;
#10;
address_ina = 24;
address_inb = 25;
data_ina = 16'h56d;
data_inb = 16'h443;
#10;
address_ina = 26;
address_inb = 27;
data_ina = 16'hfa77;
data_inb = 16'h45c;
#10;
address_ina = 28;
address_inb = 29;
data_ina = 16'hcd;
data_inb = 16'hfdf1;
#10;
address_ina = 30;
address_inb = 31;
data_ina = 16'h503;
data_inb = 16'h78;
#10;
address_ina = 32;
address_inb = 33;
data_ina = 16'h3f8;
data_inb = 16'h3fe;
#10;
address_ina = 34;
address_inb = 35;
data_ina = 16'h169;
data_inb = 16'h331;
#10;
address_ina = 36;
address_inb = 37;
data_ina = 16'h2c5;
data_inb = 16'hfd10;
#10;
address_ina = 38;
address_inb = 39;
data_ina = 16'hffab;
data_inb = 16'hfccc;
#10;
address_ina = 40;
address_inb = 41;
data_ina = 16'hfd55;
data_inb = 16'hff;
#10;
address_ina = 42;
address_inb = 43;
data_ina = 16'hfac2;
data_inb = 16'hfe27;
#10;
address_ina = 44;
address_inb = 45;
data_ina = 16'h335;
data_inb = 16'hfe03;
#10;
address_ina = 46;
address_inb = 47;
data_ina = 16'hd6;
data_inb = 16'ha1;
#10;
address_ina = 48;
address_inb = 49;
data_ina = 16'he7;
data_inb = 16'hfba0;
#10;
address_ina = 50;
address_inb = 51;
data_ina = 16'hfb6e;
data_inb = 16'h61d;
#10;
address_ina = 52;
address_inb = 53;
data_ina = 16'h347;
data_inb = 16'hfbe7;
#10;
address_ina = 54;
address_inb = 55;
data_ina = 16'hfc30;
data_inb = 16'hfc44;
#10;
address_ina = 56;
address_inb = 57;
data_ina = 16'hcd;
data_inb = 16'h62b;
#10;
address_ina = 58;
address_inb = 59;
data_ina = 16'hffa9;
data_inb = 16'hfa1d;
#10;
address_ina = 60;
address_inb = 61;
data_ina = 16'hf9d5;
data_inb = 16'hfecf;
#10;
address_ina = 62;
address_inb = 63;
data_ina = 16'hf9a6;
data_inb = 16'hff54;
#10;
address_ina = 64;
address_inb = 65;
data_ina = 16'hff1f;
data_inb = 16'h337;
#10;
address_ina = 66;
address_inb = 67;
data_ina = 16'hffe2;
data_inb = 16'h231;
#10;
address_ina = 68;
address_inb = 69;
data_ina = 16'hfe4e;
data_inb = 16'he3;
#10;
address_ina = 70;
address_inb = 71;
data_ina = 16'h5ae;
data_inb = 16'hfe3b;
#10;
address_ina = 72;
address_inb = 73;
data_ina = 16'h333;
data_inb = 16'h380;
#10;
address_ina = 74;
address_inb = 75;
data_ina = 16'h256;
data_inb = 16'hfbde;
#10;
address_ina = 76;
address_inb = 77;
data_ina = 16'hfc72;
data_inb = 16'hfa1e;
#10;
address_ina = 78;
address_inb = 79;
data_ina = 16'hfe52;
data_inb = 16'h28;
#10;
address_ina = 80;
address_inb = 81;
data_ina = 16'hfa51;
data_inb = 16'h3aa;
#10;
address_ina = 82;
address_inb = 83;
data_ina = 16'hff63;
data_inb = 16'h444;
#10;
address_ina = 84;
address_inb = 85;
data_ina = 16'hfb33;
data_inb = 16'h38c;
#10;
address_ina = 86;
address_inb = 87;
data_ina = 16'h170;
data_inb = 16'h437;
#10;
address_ina = 88;
address_inb = 89;
data_ina = 16'h32c;
data_inb = 16'hfaba;
#10;
address_ina = 90;
address_inb = 91;
data_ina = 16'hfc91;
data_inb = 16'hfe86;
#10;
address_ina = 92;
address_inb = 93;
data_ina = 16'hfea1;
data_inb = 16'h45b;
#10;
address_ina = 94;
address_inb = 95;
data_ina = 16'hfae9;
data_inb = 16'h57f;
#10;
address_ina = 96;
address_inb = 97;
data_ina = 16'hff0e;
data_inb = 16'h518;
#10;
address_ina = 98;
address_inb = 99;
data_ina = 16'h1ce;
data_inb = 16'hfbc7;
#10;
address_ina = 100;
address_inb = 101;
data_ina = 16'h1fc;
data_inb = 16'hfa05;
#10;
address_ina = 102;
address_inb = 103;
data_ina = 16'hf9f9;
data_inb = 16'h471;
#10;
address_ina = 104;
address_inb = 105;
data_ina = 16'hfff9;
data_inb = 16'hfe34;
#10;
address_ina = 106;
address_inb = 107;
data_ina = 16'h475;
data_inb = 16'hfc53;
#10;
address_ina = 108;
address_inb = 109;
data_ina = 16'hfb38;
data_inb = 16'hfbfb;
#10;
address_ina = 110;
address_inb = 111;
data_ina = 16'hfbc9;
data_inb = 16'hfb73;
#10;
address_ina = 112;
address_inb = 113;
data_ina = 16'h116;
data_inb = 16'h4d8;
#10;
address_ina = 114;
address_inb = 115;
data_ina = 16'h528;
data_inb = 16'h4a5;
#10;
address_ina = 116;
address_inb = 117;
data_ina = 16'hfbb0;
data_inb = 16'hfd55;
#10;
address_ina = 118;
address_inb = 119;
data_ina = 16'h399;
data_inb = 16'h4ff;
#10;
address_ina = 120;
address_inb = 121;
data_ina = 16'h7a;
data_inb = 16'h38f;
#10;
address_ina = 122;
address_inb = 123;
data_ina = 16'hfc50;
data_inb = 16'hff5a;
#10;
address_ina = 124;
address_inb = 125;
data_ina = 16'hf986;
data_inb = 16'h3fd;
#10;
address_ina = 126;
address_inb = 127;
data_ina = 16'h5e5;
data_inb = 16'h56f;
#10;
address_ina = 128;
address_inb = 129;
data_ina = 16'hff50;
data_inb = 16'hfbe8;
#10;
address_ina = 130;
address_inb = 131;
data_ina = 16'h166;
data_inb = 16'h305;
#10;
address_ina = 132;
address_inb = 133;
data_ina = 16'hfc9a;
data_inb = 16'h317;
#10;
address_ina = 134;
address_inb = 135;
data_ina = 16'h2c0;
data_inb = 16'hfd48;
#10;
address_ina = 136;
address_inb = 137;
data_ina = 16'h5bf;
data_inb = 16'h297;
#10;
address_ina = 138;
address_inb = 139;
data_ina = 16'h59d;
data_inb = 16'hfb63;
#10;
address_ina = 140;
address_inb = 141;
data_ina = 16'hfcf1;
data_inb = 16'h153;
#10;
address_ina = 142;
address_inb = 143;
data_ina = 16'hfefe;
data_inb = 16'h2bc;
#10;
address_ina = 144;
address_inb = 145;
data_ina = 16'h64;
data_inb = 16'hfbf3;
#10;
address_ina = 146;
address_inb = 147;
data_ina = 16'h1cc;
data_inb = 16'h294;
#10;
address_ina = 148;
address_inb = 149;
data_ina = 16'h23f;
data_inb = 16'h5f0;
#10;
address_ina = 150;
address_inb = 151;
data_ina = 16'h2ec;
data_inb = 16'hc4;
#10;
address_ina = 152;
address_inb = 153;
data_ina = 16'hd8;
data_inb = 16'heb;
#10;
address_ina = 154;
address_inb = 155;
data_ina = 16'hf985;
data_inb = 16'hffc8;
#10;
address_ina = 156;
address_inb = 157;
data_ina = 16'hff4e;
data_inb = 16'hfe23;
#10;
address_ina = 158;
address_inb = 159;
data_ina = 16'hfcc5;
data_inb = 16'hfae4;
#10;
address_ina = 160;
address_inb = 161;
data_ina = 16'hfd28;
data_inb = 16'h632;
#10;
address_ina = 162;
address_inb = 163;
data_ina = 16'h31b;
data_inb = 16'hfad7;
#10;
address_ina = 164;
address_inb = 165;
data_ina = 16'hff7d;
data_inb = 16'hfa9a;
#10;
address_ina = 166;
address_inb = 167;
data_ina = 16'h436;
data_inb = 16'hff63;
#10;
address_ina = 168;
address_inb = 169;
data_ina = 16'hfb0d;
data_inb = 16'h1a;
#10;
address_ina = 170;
address_inb = 171;
data_ina = 16'hfa97;
data_inb = 16'h648;
#10;
address_ina = 172;
address_inb = 173;
data_ina = 16'hfe77;
data_inb = 16'h1cf;
#10;
address_ina = 174;
address_inb = 175;
data_ina = 16'hff65;
data_inb = 16'h5f;
#10;
address_ina = 176;
address_inb = 177;
data_ina = 16'hff50;
data_inb = 16'h90;
#10;
address_ina = 178;
address_inb = 179;
data_ina = 16'h580;
data_inb = 16'hab;
#10;
address_ina = 180;
address_inb = 181;
data_ina = 16'h513;
data_inb = 16'h45c;
#10;
address_ina = 182;
address_inb = 183;
data_ina = 16'hfbe4;
data_inb = 16'h284;
#10;
address_ina = 184;
address_inb = 185;
data_ina = 16'h3ab;
data_inb = 16'ha4;
#10;
address_ina = 186;
address_inb = 187;
data_ina = 16'hfeac;
data_inb = 16'h3bb;
#10;
address_ina = 188;
address_inb = 189;
data_ina = 16'h435;
data_inb = 16'hfc8a;
#10;
address_ina = 190;
address_inb = 191;
data_ina = 16'hff77;
data_inb = 16'h48c;
#10;
address_ina = 192;
address_inb = 193;
data_ina = 16'hff85;
data_inb = 16'h5d5;
#10;
address_ina = 194;
address_inb = 195;
data_ina = 16'h2a4;
data_inb = 16'hfd5d;
#10;
address_ina = 196;
address_inb = 197;
data_ina = 16'h43;
data_inb = 16'hfe34;
#10;
address_ina = 198;
address_inb = 199;
data_ina = 16'hff65;
data_inb = 16'h492;
#10;
address_ina = 200;
address_inb = 201;
data_ina = 16'hfd97;
data_inb = 16'h3c4;
#10;
address_ina = 202;
address_inb = 203;
data_ina = 16'hfdeb;
data_inb = 16'h2f4;
#10;
address_ina = 204;
address_inb = 205;
data_ina = 16'h316;
data_inb = 16'hff92;
#10;
address_ina = 206;
address_inb = 207;
data_ina = 16'hfa80;
data_inb = 16'h652;
#10;
address_ina = 208;
address_inb = 209;
data_ina = 16'hfb87;
data_inb = 16'hfacd;
#10;
address_ina = 210;
address_inb = 211;
data_ina = 16'hfb95;
data_inb = 16'hfa29;
#10;
address_ina = 212;
address_inb = 213;
data_ina = 16'hfd04;
data_inb = 16'h44f;
#10;
address_ina = 214;
address_inb = 215;
data_ina = 16'h2d1;
data_inb = 16'h53d;
#10;
address_ina = 216;
address_inb = 217;
data_ina = 16'hfa05;
data_inb = 16'h4f0;
#10;
address_ina = 218;
address_inb = 219;
data_ina = 16'h28b;
data_inb = 16'hfd65;
#10;
address_ina = 220;
address_inb = 221;
data_ina = 16'h50;
data_inb = 16'h36f;
#10;
address_ina = 222;
address_inb = 223;
data_ina = 16'h30a;
data_inb = 16'h5e1;
#10;
address_ina = 224;
address_inb = 225;
data_ina = 16'ha6;
data_inb = 16'hfc6a;
#10;
address_ina = 226;
address_inb = 227;
data_ina = 16'h5ba;
data_inb = 16'h36b;
#10;
address_ina = 228;
address_inb = 229;
data_ina = 16'hff4f;
data_inb = 16'h637;
#10;
address_ina = 230;
address_inb = 231;
data_ina = 16'hfb2b;
data_inb = 16'hf986;
#10;
address_ina = 232;
address_inb = 233;
data_ina = 16'h4ef;
data_inb = 16'h1ec;
#10;
address_ina = 234;
address_inb = 235;
data_ina = 16'hf991;
data_inb = 16'hfbb3;
#10;
address_ina = 236;
address_inb = 237;
data_ina = 16'h4ed;
data_inb = 16'h556;
#10;
address_ina = 238;
address_inb = 239;
data_ina = 16'h149;
data_inb = 16'hfce0;
#10;
address_ina = 240;
address_inb = 241;
data_ina = 16'hfe4b;
data_inb = 16'hfbb7;
#10;
address_ina = 242;
address_inb = 243;
data_ina = 16'hff54;
data_inb = 16'h4a4;
#10;
address_ina = 244;
address_inb = 245;
data_ina = 16'hfc98;
data_inb = 16'h26f;
#10;
address_ina = 246;
address_inb = 247;
data_ina = 16'hff7a;
data_inb = 16'h626;
#10;
address_ina = 248;
address_inb = 249;
data_ina = 16'hfdc4;
data_inb = 16'h21a;
#10;
address_ina = 250;
address_inb = 251;
data_ina = 16'h2b9;
data_inb = 16'h5a5;
#10;
address_ina = 252;
address_inb = 253;
data_ina = 16'hfc35;
data_inb = 16'h55e;
#10;
address_ina = 254;
address_inb = 255;
data_ina = 16'h3e3;
data_inb = 16'hffea;
#10;
        wait(init_done);
        #30
        we = 0;
        // Start processing
         
		  #38000

        start = 0;



//        wait (wr_req);
//		  wait (!wr_req);
//		   rd_req = 1;
		  wait(done);
		  #20000
rd_req = 1;
        #70 
		  start = 1;
		 #80 
wait(rd_empty)
rd_req = 0;

$display("Finished the NTT test Number %d",test_num);
////Begin test number #26//////////////
rst = 1;

//#1000
start = 1;
mode = 0; //NTT 0 // INTT 1

// Reset for a few clock cycles

#1000

rst = 0;
test_num = test_num + 1;
#1000
we = 1;
address_ina = 0;
address_inb = 1;
data_ina = 16'h4c6;
data_inb = 16'ha8a;
#10;
address_ina = 2;
address_inb = 3;
data_ina = 16'h9b4;
data_inb = 16'h2ec;
#10;
address_ina = 4;
address_inb = 5;
data_ina = 16'h6f2;
data_inb = 16'h911;
#10;
address_ina = 6;
address_inb = 7;
data_ina = 16'hfa;
data_inb = 16'h7c;
#10;
address_ina = 8;
address_inb = 9;
data_ina = 16'hb1d;
data_inb = 16'h5f1;
#10;
address_ina = 10;
address_inb = 11;
data_ina = 16'h2bb;
data_inb = 16'h388;
#10;
address_ina = 12;
address_inb = 13;
data_ina = 16'h4fa;
data_inb = 16'h16c;
#10;
address_ina = 14;
address_inb = 15;
data_ina = 16'h6d2;
data_inb = 16'h778;
#10;
address_ina = 16;
address_inb = 17;
data_ina = 16'hc00;
data_inb = 16'h899;
#10;
address_ina = 18;
address_inb = 19;
data_ina = 16'h4ac;
data_inb = 16'h39f;
#10;
address_ina = 20;
address_inb = 21;
data_ina = 16'hbb9;
data_inb = 16'h87f;
#10;
address_ina = 22;
address_inb = 23;
data_ina = 16'h6c5;
data_inb = 16'h1d4;
#10;
address_ina = 24;
address_inb = 25;
data_ina = 16'hced;
data_inb = 16'h2d2;
#10;
address_ina = 26;
address_inb = 27;
data_ina = 16'h8b0;
data_inb = 16'h673;
#10;
address_ina = 28;
address_inb = 29;
data_ina = 16'h5b4;
data_inb = 16'h660;
#10;
address_ina = 30;
address_inb = 31;
data_ina = 16'h39b;
data_inb = 16'h385;
#10;
address_ina = 32;
address_inb = 33;
data_ina = 16'h62;
data_inb = 16'h462;
#10;
address_ina = 34;
address_inb = 35;
data_ina = 16'h6b;
data_inb = 16'h72a;
#10;
address_ina = 36;
address_inb = 37;
data_ina = 16'h625;
data_inb = 16'h179;
#10;
address_ina = 38;
address_inb = 39;
data_ina = 16'h52e;
data_inb = 16'h4cd;
#10;
address_ina = 40;
address_inb = 41;
data_ina = 16'hc27;
data_inb = 16'h0;
#10;
address_ina = 42;
address_inb = 43;
data_ina = 16'haf2;
data_inb = 16'h347;
#10;
address_ina = 44;
address_inb = 45;
data_ina = 16'he0;
data_inb = 16'h579;
#10;
address_ina = 46;
address_inb = 47;
data_ina = 16'ha9b;
data_inb = 16'hcf7;
#10;
address_ina = 48;
address_inb = 49;
data_ina = 16'h7c9;
data_inb = 16'h354;
#10;
address_ina = 50;
address_inb = 51;
data_ina = 16'hcea;
data_inb = 16'h9d1;
#10;
address_ina = 52;
address_inb = 53;
data_ina = 16'h12e;
data_inb = 16'h3e0;
#10;
address_ina = 54;
address_inb = 55;
data_ina = 16'hcc3;
data_inb = 16'h8e4;
#10;
address_ina = 56;
address_inb = 57;
data_ina = 16'h7;
data_inb = 16'h38e;
#10;
address_ina = 58;
address_inb = 59;
data_ina = 16'ha1c;
data_inb = 16'h320;
#10;
address_ina = 60;
address_inb = 61;
data_ina = 16'h5de;
data_inb = 16'h9ce;
#10;
address_ina = 62;
address_inb = 63;
data_ina = 16'h670;
data_inb = 16'h6d8;
#10;
address_ina = 64;
address_inb = 65;
data_ina = 16'h26d;
data_inb = 16'h84e;
#10;
address_ina = 66;
address_inb = 67;
data_ina = 16'h57c;
data_inb = 16'h785;
#10;
address_ina = 68;
address_inb = 69;
data_ina = 16'h38e;
data_inb = 16'hab1;
#10;
address_ina = 70;
address_inb = 71;
data_ina = 16'h6fc;
data_inb = 16'ha1c;
#10;
address_ina = 72;
address_inb = 73;
data_ina = 16'h159;
data_inb = 16'hcdd;
#10;
address_ina = 74;
address_inb = 75;
data_ina = 16'h983;
data_inb = 16'h1ee;
#10;
address_ina = 76;
address_inb = 77;
data_ina = 16'hb16;
data_inb = 16'h4bd;
#10;
address_ina = 78;
address_inb = 79;
data_ina = 16'h650;
data_inb = 16'h5b;
#10;
address_ina = 80;
address_inb = 81;
data_ina = 16'h504;
data_inb = 16'ha74;
#10;
address_ina = 82;
address_inb = 83;
data_ina = 16'h35e;
data_inb = 16'hbb5;
#10;
address_ina = 84;
address_inb = 85;
data_ina = 16'h81a;
data_inb = 16'h2ce;
#10;
address_ina = 86;
address_inb = 87;
data_ina = 16'h716;
data_inb = 16'h7ac;
#10;
address_ina = 88;
address_inb = 89;
data_ina = 16'hbaf;
data_inb = 16'h622;
#10;
address_ina = 90;
address_inb = 91;
data_ina = 16'h882;
data_inb = 16'haab;
#10;
address_ina = 92;
address_inb = 93;
data_ina = 16'h97c;
data_inb = 16'h4ea;
#10;
address_ina = 94;
address_inb = 95;
data_ina = 16'h86f;
data_inb = 16'h65d;
#10;
address_ina = 96;
address_inb = 97;
data_ina = 16'h73d;
data_inb = 16'h948;
#10;
address_ina = 98;
address_inb = 99;
data_ina = 16'h61c;
data_inb = 16'h733;
#10;
address_ina = 100;
address_inb = 101;
data_ina = 16'h8cd;
data_inb = 16'h155;
#10;
address_ina = 102;
address_inb = 103;
data_ina = 16'hc5b;
data_inb = 16'hb57;
#10;
address_ina = 104;
address_inb = 105;
data_ina = 16'h44;
data_inb = 16'h824;
#10;
address_ina = 106;
address_inb = 107;
data_ina = 16'h615;
data_inb = 16'h85e;
#10;
address_ina = 108;
address_inb = 109;
data_ina = 16'h781;
data_inb = 16'h17;
#10;
address_ina = 110;
address_inb = 111;
data_ina = 16'h2c1;
data_inb = 16'h302;
#10;
address_ina = 112;
address_inb = 113;
data_ina = 16'h2ce;
data_inb = 16'hb5a;
#10;
address_ina = 114;
address_inb = 115;
data_ina = 16'ha02;
data_inb = 16'hbe6;
#10;
address_ina = 116;
address_inb = 117;
data_ina = 16'hcea;
data_inb = 16'hc5b;
#10;
address_ina = 118;
address_inb = 119;
data_ina = 16'h719;
data_inb = 16'h77b;
#10;
address_ina = 120;
address_inb = 121;
data_ina = 16'h189;
data_inb = 16'hb0;
#10;
address_ina = 122;
address_inb = 123;
data_ina = 16'hc92;
data_inb = 16'hc7f;
#10;
address_ina = 124;
address_inb = 125;
data_ina = 16'hb3d;
data_inb = 16'h294;
#10;
address_ina = 126;
address_inb = 127;
data_ina = 16'ha1c;
data_inb = 16'h93f;
#10;
address_ina = 128;
address_inb = 129;
data_ina = 16'h15f;
data_inb = 16'ha2c;
#10;
address_ina = 130;
address_inb = 131;
data_ina = 16'h21f;
data_inb = 16'h7c9;
#10;
address_ina = 132;
address_inb = 133;
data_ina = 16'hc34;
data_inb = 16'h451;
#10;
address_ina = 134;
address_inb = 135;
data_ina = 16'h81a;
data_inb = 16'hc9f;
#10;
address_ina = 136;
address_inb = 137;
data_ina = 16'ha5a;
data_inb = 16'h148;
#10;
address_ina = 138;
address_inb = 139;
data_ina = 16'hc62;
data_inb = 16'h111;
#10;
address_ina = 140;
address_inb = 141;
data_ina = 16'hc8c;
data_inb = 16'h899;
#10;
address_ina = 142;
address_inb = 143;
data_ina = 16'h586;
data_inb = 16'h764;
#10;
address_ina = 144;
address_inb = 145;
data_ina = 16'h410;
data_inb = 16'h862;
#10;
address_ina = 146;
address_inb = 147;
data_ina = 16'h1bd;
data_inb = 16'h921;
#10;
address_ina = 148;
address_inb = 149;
data_ina = 16'hce4;
data_inb = 16'h395;
#10;
address_ina = 150;
address_inb = 151;
data_ina = 16'h229;
data_inb = 16'h458;
#10;
address_ina = 152;
address_inb = 153;
data_ina = 16'hc51;
data_inb = 16'h848;
#10;
address_ina = 154;
address_inb = 155;
data_ina = 16'h62f;
data_inb = 16'h91e;
#10;
address_ina = 156;
address_inb = 157;
data_ina = 16'h697;
data_inb = 16'h942;
#10;
address_ina = 158;
address_inb = 159;
data_ina = 16'h7;
data_inb = 16'h44e;
#10;
address_ina = 160;
address_inb = 161;
data_ina = 16'h3b2;
data_inb = 16'hc48;
#10;
address_ina = 162;
address_inb = 163;
data_ina = 16'h862;
data_inb = 16'h521;
#10;
address_ina = 164;
address_inb = 165;
data_ina = 16'h7b9;
data_inb = 16'h9a7;
#10;
address_ina = 166;
address_inb = 167;
data_ina = 16'h694;
data_inb = 16'h4e;
#10;
address_ina = 168;
address_inb = 169;
data_ina = 16'h632;
data_inb = 16'h625;
#10;
address_ina = 170;
address_inb = 171;
data_ina = 16'h6dc;
data_inb = 16'h8e4;
#10;
address_ina = 172;
address_inb = 173;
data_ina = 16'hb81;
data_inb = 16'h11e;
#10;
address_ina = 174;
address_inb = 175;
data_ina = 16'h114;
data_inb = 16'h4f1;
#10;
address_ina = 176;
address_inb = 177;
data_ina = 16'h4fa;
data_inb = 16'h280;
#10;
address_ina = 178;
address_inb = 179;
data_ina = 16'hce4;
data_inb = 16'h8c6;
#10;
address_ina = 180;
address_inb = 181;
data_ina = 16'h3dc;
data_inb = 16'h5b0;
#10;
address_ina = 182;
address_inb = 183;
data_ina = 16'h54c;
data_inb = 16'h44b;
#10;
address_ina = 184;
address_inb = 185;
data_ina = 16'h7ed;
data_inb = 16'h625;
#10;
address_ina = 186;
address_inb = 187;
data_ina = 16'h6b5;
data_inb = 16'hb2a;
#10;
address_ina = 188;
address_inb = 189;
data_ina = 16'h4c6;
data_inb = 16'h673;
#10;
address_ina = 190;
address_inb = 191;
data_ina = 16'hba2;
data_inb = 16'h478;
#10;
address_ina = 192;
address_inb = 193;
data_ina = 16'h176;
data_inb = 16'h8ea;
#10;
address_ina = 194;
address_inb = 195;
data_ina = 16'hbb2;
data_inb = 16'h7ac;
#10;
address_ina = 196;
address_inb = 197;
data_ina = 16'ha43;
data_inb = 16'h351;
#10;
address_ina = 198;
address_inb = 199;
data_ina = 16'h68;
data_inb = 16'hcdd;
#10;
address_ina = 200;
address_inb = 201;
data_ina = 16'h67d;
data_inb = 16'hc82;
#10;
address_ina = 202;
address_inb = 203;
data_ina = 16'h3ed;
data_inb = 16'hb9;
#10;
address_ina = 204;
address_inb = 205;
data_ina = 16'h747;
data_inb = 16'hb64;
#10;
address_ina = 206;
address_inb = 207;
data_ina = 16'hb67;
data_inb = 16'hc0a;
#10;
address_ina = 208;
address_inb = 209;
data_ina = 16'h12b;
data_inb = 16'h559;
#10;
address_ina = 210;
address_inb = 211;
data_ina = 16'h482;
data_inb = 16'h23f;
#10;
address_ina = 212;
address_inb = 213;
data_ina = 16'h33a;
data_inb = 16'hc5b;
#10;
address_ina = 214;
address_inb = 215;
data_ina = 16'h6d5;
data_inb = 16'h7f0;
#10;
address_ina = 216;
address_inb = 217;
data_ina = 16'h183;
data_inb = 16'h6ff;
#10;
address_ina = 218;
address_inb = 219;
data_ina = 16'hcb9;
data_inb = 16'habb;
#10;
address_ina = 220;
address_inb = 221;
data_ina = 16'h1d4;
data_inb = 16'h10e;
#10;
address_ina = 222;
address_inb = 223;
data_ina = 16'h3f0;
data_inb = 16'hc2e;
#10;
address_ina = 224;
address_inb = 225;
data_ina = 16'hb78;
data_inb = 16'h84e;
#10;
address_ina = 226;
address_inb = 227;
data_ina = 16'hda;
data_inb = 16'ha84;
#10;
address_ina = 228;
address_inb = 229;
data_ina = 16'h55c;
data_inb = 16'h841;
#10;
address_ina = 230;
address_inb = 231;
data_ina = 16'h77e;
data_inb = 16'h7fa;
#10;
address_ina = 232;
address_inb = 233;
data_ina = 16'h74d;
data_inb = 16'hb9f;
#10;
address_ina = 234;
address_inb = 235;
data_ina = 16'ha26;
data_inb = 16'h9db;
#10;
address_ina = 236;
address_inb = 237;
data_ina = 16'hb4d;
data_inb = 16'h25d;
#10;
address_ina = 238;
address_inb = 239;
data_ina = 16'h40d;
data_inb = 16'h629;
#10;
address_ina = 240;
address_inb = 241;
data_ina = 16'h938;
data_inb = 16'h800;
#10;
address_ina = 242;
address_inb = 243;
data_ina = 16'h649;
data_inb = 16'h3f3;
#10;
address_ina = 244;
address_inb = 245;
data_ina = 16'h72d;
data_inb = 16'h1ba;
#10;
address_ina = 246;
address_inb = 247;
data_ina = 16'hac;
data_inb = 16'h4b0;
#10;
address_ina = 248;
address_inb = 249;
data_ina = 16'h169;
data_inb = 16'h580;
#10;
address_ina = 250;
address_inb = 251;
data_ina = 16'h43e;
data_inb = 16'h681;
#10;
address_ina = 252;
address_inb = 253;
data_ina = 16'h56f;
data_inb = 16'h4b3;
#10;
address_ina = 254;
address_inb = 255;
data_ina = 16'h95f;
data_inb = 16'h24c;
#10;
        wait(init_done);
        #30
        we = 0;
        // Start processing
         
		  #38000

        start = 0;



//        wait (wr_req);
//		  wait (!wr_req);
//		   rd_req = 1;
		  wait(done);
		  #20000
rd_req = 1;
        #70 
		  start = 1;
		 #80 
wait(rd_empty)
rd_req = 0;

$display("Finished the NTT test Number %d",test_num);
////Begin test number #27//////////////
rst = 1;

//#1000
start = 1;
mode = 0; //NTT 0 // INTT 1

// Reset for a few clock cycles

#1000

rst = 0;
test_num = test_num + 1;
#1000
we = 1;
address_ina = 0;
address_inb = 1;
data_ina = 16'hb2a;
data_inb = 16'h2a7;
#10;
address_ina = 2;
address_inb = 3;
data_ina = 16'h1d1;
data_inb = 16'h132;
#10;
address_ina = 4;
address_inb = 5;
data_ina = 16'hb3d;
data_inb = 16'h36b;
#10;
address_ina = 6;
address_inb = 7;
data_ina = 16'h6c2;
data_inb = 16'h892;
#10;
address_ina = 8;
address_inb = 9;
data_ina = 16'h9f5;
data_inb = 16'h333;
#10;
address_ina = 10;
address_inb = 11;
data_ina = 16'h3dc;
data_inb = 16'h663;
#10;
address_ina = 12;
address_inb = 13;
data_ina = 16'hc0;
data_inb = 16'h62;
#10;
address_ina = 14;
address_inb = 15;
data_ina = 16'h14;
data_inb = 16'h1a;
#10;
address_ina = 16;
address_inb = 17;
data_ina = 16'hb61;
data_inb = 16'h489;
#10;
address_ina = 18;
address_inb = 19;
data_ina = 16'h3b9;
data_inb = 16'h59a;
#10;
address_ina = 20;
address_inb = 21;
data_ina = 16'h27;
data_inb = 16'hced;
#10;
address_ina = 22;
address_inb = 23;
data_ina = 16'h24;
data_inb = 16'habb;
#10;
address_ina = 24;
address_inb = 25;
data_ina = 16'h364;
data_inb = 16'hbf6;
#10;
address_ina = 26;
address_inb = 27;
data_ina = 16'h792;
data_inb = 16'hbac;
#10;
address_ina = 28;
address_inb = 29;
data_ina = 16'hfe;
data_inb = 16'h18d;
#10;
address_ina = 30;
address_inb = 31;
data_ina = 16'h8fe;
data_inb = 16'h6ff;
#10;
address_ina = 32;
address_inb = 33;
data_ina = 16'h7ac;
data_inb = 16'h952;
#10;
address_ina = 34;
address_inb = 35;
data_ina = 16'h93f;
data_inb = 16'ha;
#10;
address_ina = 36;
address_inb = 37;
data_ina = 16'h5de;
data_inb = 16'h29a;
#10;
address_ina = 38;
address_inb = 39;
data_ina = 16'hc44;
data_inb = 16'h72;
#10;
address_ina = 40;
address_inb = 41;
data_ina = 16'h4f4;
data_inb = 16'h48c;
#10;
address_ina = 42;
address_inb = 43;
data_ina = 16'h1c7;
data_inb = 16'h215;
#10;
address_ina = 44;
address_inb = 45;
data_ina = 16'h4e0;
data_inb = 16'h98d;
#10;
address_ina = 46;
address_inb = 47;
data_ina = 16'h8b0;
data_inb = 16'ha5a;
#10;
address_ina = 48;
address_inb = 49;
data_ina = 16'had2;
data_inb = 16'h928;
#10;
address_ina = 50;
address_inb = 51;
data_ina = 16'h400;
data_inb = 16'h12b;
#10;
address_ina = 52;
address_inb = 53;
data_ina = 16'h1fe;
data_inb = 16'h9c1;
#10;
address_ina = 54;
address_inb = 55;
data_ina = 16'h385;
data_inb = 16'h280;
#10;
address_ina = 56;
address_inb = 57;
data_ina = 16'h740;
data_inb = 16'hba8;
#10;
address_ina = 58;
address_inb = 59;
data_ina = 16'h434;
data_inb = 16'h14c;
#10;
address_ina = 60;
address_inb = 61;
data_ina = 16'hb2d;
data_inb = 16'h2d5;
#10;
address_ina = 62;
address_inb = 63;
data_ina = 16'hcc0;
data_inb = 16'h2e8;
#10;
address_ina = 64;
address_inb = 65;
data_ina = 16'hbb2;
data_inb = 16'h9a7;
#10;
address_ina = 66;
address_inb = 67;
data_ina = 16'h5d7;
data_inb = 16'h62f;
#10;
address_ina = 68;
address_inb = 69;
data_ina = 16'h3e0;
data_inb = 16'h684;
#10;
address_ina = 70;
address_inb = 71;
data_ina = 16'h969;
data_inb = 16'h2d8;
#10;
address_ina = 72;
address_inb = 73;
data_ina = 16'h566;
data_inb = 16'h49c;
#10;
address_ina = 74;
address_inb = 75;
data_ina = 16'h250;
data_inb = 16'h4d7;
#10;
address_ina = 76;
address_inb = 77;
data_ina = 16'h75a;
data_inb = 16'ha70;
#10;
address_ina = 78;
address_inb = 79;
data_ina = 16'h5a0;
data_inb = 16'h6a4;
#10;
address_ina = 80;
address_inb = 81;
data_ina = 16'hb1d;
data_inb = 16'h19a;
#10;
address_ina = 82;
address_inb = 83;
data_ina = 16'he4;
data_inb = 16'h932;
#10;
address_ina = 84;
address_inb = 85;
data_ina = 16'h5fe;
data_inb = 16'hbe3;
#10;
address_ina = 86;
address_inb = 87;
data_ina = 16'hcfe;
data_inb = 16'hb1d;
#10;
address_ina = 88;
address_inb = 89;
data_ina = 16'h87f;
data_inb = 16'h5a7;
#10;
address_ina = 90;
address_inb = 91;
data_ina = 16'ha40;
data_inb = 16'hcfa;
#10;
address_ina = 92;
address_inb = 93;
data_ina = 16'haa1;
data_inb = 16'hb5a;
#10;
address_ina = 94;
address_inb = 95;
data_ina = 16'h6fc;
data_inb = 16'h889;
#10;
address_ina = 96;
address_inb = 97;
data_ina = 16'h96;
data_inb = 16'haa4;
#10;
address_ina = 98;
address_inb = 99;
data_ina = 16'h44b;
data_inb = 16'hfe;
#10;
address_ina = 100;
address_inb = 101;
data_ina = 16'h2a;
data_inb = 16'h3c9;
#10;
address_ina = 102;
address_inb = 103;
data_ina = 16'h7a2;
data_inb = 16'h3d9;
#10;
address_ina = 104;
address_inb = 105;
data_ina = 16'h9a3;
data_inb = 16'h3bc;
#10;
address_ina = 106;
address_inb = 107;
data_ina = 16'hced;
data_inb = 16'h2cb;
#10;
address_ina = 108;
address_inb = 109;
data_ina = 16'ha91;
data_inb = 16'h84e;
#10;
address_ina = 110;
address_inb = 111;
data_ina = 16'h5e;
data_inb = 16'h56c;
#10;
address_ina = 112;
address_inb = 113;
data_ina = 16'h3b9;
data_inb = 16'h778;
#10;
address_ina = 114;
address_inb = 115;
data_ina = 16'hc1a;
data_inb = 16'h88f;
#10;
address_ina = 116;
address_inb = 117;
data_ina = 16'h1ca;
data_inb = 16'hc0;
#10;
address_ina = 118;
address_inb = 119;
data_ina = 16'h6bb;
data_inb = 16'h52e;
#10;
address_ina = 120;
address_inb = 121;
data_ina = 16'h788;
data_inb = 16'h1f5;
#10;
address_ina = 122;
address_inb = 123;
data_ina = 16'hb9f;
data_inb = 16'h51b;
#10;
address_ina = 124;
address_inb = 125;
data_ina = 16'h378;
data_inb = 16'hafc;
#10;
address_ina = 126;
address_inb = 127;
data_ina = 16'ha33;
data_inb = 16'h329;
#10;
address_ina = 128;
address_inb = 129;
data_ina = 16'h263;
data_inb = 16'hf1;
#10;
address_ina = 130;
address_inb = 131;
data_ina = 16'h90e;
data_inb = 16'h34a;
#10;
address_ina = 132;
address_inb = 133;
data_ina = 16'h69b;
data_inb = 16'h6bb;
#10;
address_ina = 134;
address_inb = 135;
data_ina = 16'h87c;
data_inb = 16'h2c8;
#10;
address_ina = 136;
address_inb = 137;
data_ina = 16'hbf6;
data_inb = 16'h8e0;
#10;
address_ina = 138;
address_inb = 139;
data_ina = 16'h92e;
data_inb = 16'h7c;
#10;
address_ina = 140;
address_inb = 141;
data_ina = 16'h7c;
data_inb = 16'h218;
#10;
address_ina = 142;
address_inb = 143;
data_ina = 16'h208;
data_inb = 16'h643;
#10;
address_ina = 144;
address_inb = 145;
data_ina = 16'h8e4;
data_inb = 16'h7c6;
#10;
address_ina = 146;
address_inb = 147;
data_ina = 16'hca9;
data_inb = 16'h1f8;
#10;
address_ina = 148;
address_inb = 149;
data_ina = 16'h472;
data_inb = 16'h9db;
#10;
address_ina = 150;
address_inb = 151;
data_ina = 16'ha6d;
data_inb = 16'hbf6;
#10;
address_ina = 152;
address_inb = 153;
data_ina = 16'h7fd;
data_inb = 16'h69e;
#10;
address_ina = 154;
address_inb = 155;
data_ina = 16'h3c9;
data_inb = 16'h82a;
#10;
address_ina = 156;
address_inb = 157;
data_ina = 16'h959;
data_inb = 16'h472;
#10;
address_ina = 158;
address_inb = 159;
data_ina = 16'h1b0;
data_inb = 16'h3af;
#10;
address_ina = 160;
address_inb = 161;
data_ina = 16'h8f1;
data_inb = 16'h33d;
#10;
address_ina = 162;
address_inb = 163;
data_ina = 16'h31;
data_inb = 16'hb9;
#10;
address_ina = 164;
address_inb = 165;
data_ina = 16'hbe3;
data_inb = 16'h340;
#10;
address_ina = 166;
address_inb = 167;
data_ina = 16'h31;
data_inb = 16'h270;
#10;
address_ina = 168;
address_inb = 169;
data_ina = 16'h751;
data_inb = 16'hb10;
#10;
address_ina = 170;
address_inb = 171;
data_ina = 16'hb7e;
data_inb = 16'h87c;
#10;
address_ina = 172;
address_inb = 173;
data_ina = 16'h7c2;
data_inb = 16'h7d9;
#10;
address_ina = 174;
address_inb = 175;
data_ina = 16'h6d5;
data_inb = 16'h36b;
#10;
address_ina = 176;
address_inb = 177;
data_ina = 16'hc7f;
data_inb = 16'h138;
#10;
address_ina = 178;
address_inb = 179;
data_ina = 16'h93f;
data_inb = 16'h72a;
#10;
address_ina = 180;
address_inb = 181;
data_ina = 16'habe;
data_inb = 16'h4ed;
#10;
address_ina = 182;
address_inb = 183;
data_ina = 16'hc17;
data_inb = 16'h9a7;
#10;
address_ina = 184;
address_inb = 185;
data_ina = 16'h659;
data_inb = 16'had5;
#10;
address_ina = 186;
address_inb = 187;
data_ina = 16'h1d7;
data_inb = 16'h183;
#10;
address_ina = 188;
address_inb = 189;
data_ina = 16'hc4e;
data_inb = 16'h13b;
#10;
address_ina = 190;
address_inb = 191;
data_ina = 16'h2e2;
data_inb = 16'hc8c;
#10;
address_ina = 192;
address_inb = 193;
data_ina = 16'h319;
data_inb = 16'haa1;
#10;
address_ina = 194;
address_inb = 195;
data_ina = 16'h34a;
data_inb = 16'h367;
#10;
address_ina = 196;
address_inb = 197;
data_ina = 16'hb5e;
data_inb = 16'h2fc;
#10;
address_ina = 198;
address_inb = 199;
data_ina = 16'h7cc;
data_inb = 16'h9b0;
#10;
address_ina = 200;
address_inb = 201;
data_ina = 16'h72a;
data_inb = 16'h6f;
#10;
address_ina = 202;
address_inb = 203;
data_ina = 16'hab5;
data_inb = 16'h7ac;
#10;
address_ina = 204;
address_inb = 205;
data_ina = 16'h0;
data_inb = 16'hc68;
#10;
address_ina = 206;
address_inb = 207;
data_ina = 16'h104;
data_inb = 16'h535;
#10;
address_ina = 208;
address_inb = 209;
data_ina = 16'h35e;
data_inb = 16'h8a3;
#10;
address_ina = 210;
address_inb = 211;
data_ina = 16'h28d;
data_inb = 16'hba8;
#10;
address_ina = 212;
address_inb = 213;
data_ina = 16'hced;
data_inb = 16'h66a;
#10;
address_ina = 214;
address_inb = 215;
data_ina = 16'h5f8;
data_inb = 16'hb7b;
#10;
address_ina = 216;
address_inb = 217;
data_ina = 16'h837;
data_inb = 16'h8dd;
#10;
address_ina = 218;
address_inb = 219;
data_ina = 16'h9c7;
data_inb = 16'h9b4;
#10;
address_ina = 220;
address_inb = 221;
data_ina = 16'h521;
data_inb = 16'hcd0;
#10;
address_ina = 222;
address_inb = 223;
data_ina = 16'h6e5;
data_inb = 16'h566;
#10;
address_ina = 224;
address_inb = 225;
data_ina = 16'hc1a;
data_inb = 16'hb6e;
#10;
address_ina = 226;
address_inb = 227;
data_ina = 16'h51e;
data_inb = 16'he0;
#10;
address_ina = 228;
address_inb = 229;
data_ina = 16'h3dc;
data_inb = 16'h914;
#10;
address_ina = 230;
address_inb = 231;
data_ina = 16'h2c1;
data_inb = 16'h26a;
#10;
address_ina = 232;
address_inb = 233;
data_ina = 16'h76b;
data_inb = 16'h91e;
#10;
address_ina = 234;
address_inb = 235;
data_ina = 16'h7fa;
data_inb = 16'h7fa;
#10;
address_ina = 236;
address_inb = 237;
data_ina = 16'hcb0;
data_inb = 16'h90e;
#10;
address_ina = 238;
address_inb = 239;
data_ina = 16'h41d;
data_inb = 16'h687;
#10;
address_ina = 240;
address_inb = 241;
data_ina = 16'h99d;
data_inb = 16'h180;
#10;
address_ina = 242;
address_inb = 243;
data_ina = 16'h966;
data_inb = 16'hc3e;
#10;
address_ina = 244;
address_inb = 245;
data_ina = 16'h993;
data_inb = 16'h1d1;
#10;
address_ina = 246;
address_inb = 247;
data_ina = 16'h482;
data_inb = 16'h2bb;
#10;
address_ina = 248;
address_inb = 249;
data_ina = 16'hba2;
data_inb = 16'h43b;
#10;
address_ina = 250;
address_inb = 251;
data_ina = 16'h9fb;
data_inb = 16'hadc;
#10;
address_ina = 252;
address_inb = 253;
data_ina = 16'h1ba;
data_inb = 16'h72d;
#10;
address_ina = 254;
address_inb = 255;
data_ina = 16'h827;
data_inb = 16'h8bd;
#10;
        wait(init_done);
        #30
        we = 0;
        // Start processing
         
		  #38000

        start = 0;



//        wait (wr_req);
//		  wait (!wr_req);
//		   rd_req = 1;
		  wait(done);
		  #20000
rd_req = 1;
        #70 
		  start = 1;
		 #80 
wait(rd_empty)
rd_req = 0;

$display("Finished the NTT test Number %d",test_num);
////Begin test number #28//////////////
rst = 1;

//#1000
start = 1;
mode = 1; //NTT 0 // INTT 1

// Reset for a few clock cycles

#1000

rst = 0;
test_num = test_num + 1;
#1000
we = 1;
address_ina = 0;
address_inb = 1;
data_ina = 16'h4c;
data_inb = 16'hfe96;
#10;
address_ina = 2;
address_inb = 3;
data_ina = 16'h3e4;
data_inb = 16'h299;
#10;
address_ina = 4;
address_inb = 5;
data_ina = 16'h4aa;
data_inb = 16'hfc9c;
#10;
address_ina = 6;
address_inb = 7;
data_ina = 16'h550;
data_inb = 16'h50e;
#10;
address_ina = 8;
address_inb = 9;
data_ina = 16'h210;
data_inb = 16'h1c4;
#10;
address_ina = 10;
address_inb = 11;
data_ina = 16'hfc4f;
data_inb = 16'hfcd3;
#10;
address_ina = 12;
address_inb = 13;
data_ina = 16'hfd14;
data_inb = 16'hfa2b;
#10;
address_ina = 14;
address_inb = 15;
data_ina = 16'h3ac;
data_inb = 16'h60b;
#10;
address_ina = 16;
address_inb = 17;
data_ina = 16'h3c3;
data_inb = 16'hff3d;
#10;
address_ina = 18;
address_inb = 19;
data_ina = 16'h69;
data_inb = 16'h65b;
#10;
address_ina = 20;
address_inb = 21;
data_ina = 16'hfe7a;
data_inb = 16'hff3c;
#10;
address_ina = 22;
address_inb = 23;
data_ina = 16'h3c6;
data_inb = 16'hf9d8;
#10;
address_ina = 24;
address_inb = 25;
data_ina = 16'hff4f;
data_inb = 16'hfe67;
#10;
address_ina = 26;
address_inb = 27;
data_ina = 16'hfdb4;
data_inb = 16'h442;
#10;
address_ina = 28;
address_inb = 29;
data_ina = 16'h517;
data_inb = 16'hfff3;
#10;
address_ina = 30;
address_inb = 31;
data_ina = 16'h35f;
data_inb = 16'h621;
#10;
address_ina = 32;
address_inb = 33;
data_ina = 16'hf984;
data_inb = 16'hfd5d;
#10;
address_ina = 34;
address_inb = 35;
data_ina = 16'h50d;
data_inb = 16'hfcc8;
#10;
address_ina = 36;
address_inb = 37;
data_ina = 16'hff99;
data_inb = 16'h512;
#10;
address_ina = 38;
address_inb = 39;
data_ina = 16'h4b;
data_inb = 16'h342;
#10;
address_ina = 40;
address_inb = 41;
data_ina = 16'h458;
data_inb = 16'hfdc7;
#10;
address_ina = 42;
address_inb = 43;
data_ina = 16'hfdd3;
data_inb = 16'hfeb5;
#10;
address_ina = 44;
address_inb = 45;
data_ina = 16'h189;
data_inb = 16'hfe64;
#10;
address_ina = 46;
address_inb = 47;
data_ina = 16'h20;
data_inb = 16'hfa97;
#10;
address_ina = 48;
address_inb = 49;
data_ina = 16'h43c;
data_inb = 16'h41e;
#10;
address_ina = 50;
address_inb = 51;
data_ina = 16'hfb0d;
data_inb = 16'h679;
#10;
address_ina = 52;
address_inb = 53;
data_ina = 16'h3a5;
data_inb = 16'h2d1;
#10;
address_ina = 54;
address_inb = 55;
data_ina = 16'hfc04;
data_inb = 16'h42e;
#10;
address_ina = 56;
address_inb = 57;
data_ina = 16'h534;
data_inb = 16'hfc6a;
#10;
address_ina = 58;
address_inb = 59;
data_ina = 16'h5f8;
data_inb = 16'h426;
#10;
address_ina = 60;
address_inb = 61;
data_ina = 16'h404;
data_inb = 16'hfc21;
#10;
address_ina = 62;
address_inb = 63;
data_ina = 16'h1b1;
data_inb = 16'h2af;
#10;
address_ina = 64;
address_inb = 65;
data_ina = 16'hfe23;
data_inb = 16'h46d;
#10;
address_ina = 66;
address_inb = 67;
data_ina = 16'hfa7d;
data_inb = 16'hff19;
#10;
address_ina = 68;
address_inb = 69;
data_ina = 16'hfab1;
data_inb = 16'h3c7;
#10;
address_ina = 70;
address_inb = 71;
data_ina = 16'h1da;
data_inb = 16'hfa38;
#10;
address_ina = 72;
address_inb = 73;
data_ina = 16'hface;
data_inb = 16'h123;
#10;
address_ina = 74;
address_inb = 75;
data_ina = 16'h5ff;
data_inb = 16'hfa3b;
#10;
address_ina = 76;
address_inb = 77;
data_ina = 16'hfef6;
data_inb = 16'hfdaf;
#10;
address_ina = 78;
address_inb = 79;
data_ina = 16'hff68;
data_inb = 16'hffe7;
#10;
address_ina = 80;
address_inb = 81;
data_ina = 16'hfcc7;
data_inb = 16'h24;
#10;
address_ina = 82;
address_inb = 83;
data_ina = 16'h3e2;
data_inb = 16'hfd95;
#10;
address_ina = 84;
address_inb = 85;
data_ina = 16'h303;
data_inb = 16'hfa63;
#10;
address_ina = 86;
address_inb = 87;
data_ina = 16'h8e;
data_inb = 16'hfbd1;
#10;
address_ina = 88;
address_inb = 89;
data_ina = 16'hfc67;
data_inb = 16'hfaa8;
#10;
address_ina = 90;
address_inb = 91;
data_ina = 16'hfb61;
data_inb = 16'hfd77;
#10;
address_ina = 92;
address_inb = 93;
data_ina = 16'hfaf2;
data_inb = 16'h50d;
#10;
address_ina = 94;
address_inb = 95;
data_ina = 16'hfed4;
data_inb = 16'hfa26;
#10;
address_ina = 96;
address_inb = 97;
data_ina = 16'hffdc;
data_inb = 16'hfdc9;
#10;
address_ina = 98;
address_inb = 99;
data_ina = 16'h4c1;
data_inb = 16'hfe7f;
#10;
address_ina = 100;
address_inb = 101;
data_ina = 16'h677;
data_inb = 16'hfb4e;
#10;
address_ina = 102;
address_inb = 103;
data_ina = 16'hfdd1;
data_inb = 16'h168;
#10;
address_ina = 104;
address_inb = 105;
data_ina = 16'hfc46;
data_inb = 16'hfd28;
#10;
address_ina = 106;
address_inb = 107;
data_ina = 16'hfb1c;
data_inb = 16'h5cb;
#10;
address_ina = 108;
address_inb = 109;
data_ina = 16'hfc7b;
data_inb = 16'h2f7;
#10;
address_ina = 110;
address_inb = 111;
data_ina = 16'hfdcc;
data_inb = 16'hfb85;
#10;
address_ina = 112;
address_inb = 113;
data_ina = 16'h3d9;
data_inb = 16'h115;
#10;
address_ina = 114;
address_inb = 115;
data_ina = 16'h327;
data_inb = 16'hfdb4;
#10;
address_ina = 116;
address_inb = 117;
data_ina = 16'hfe0f;
data_inb = 16'h59b;
#10;
address_ina = 118;
address_inb = 119;
data_ina = 16'h477;
data_inb = 16'hffbc;
#10;
address_ina = 120;
address_inb = 121;
data_ina = 16'h61d;
data_inb = 16'hfb4d;
#10;
address_ina = 122;
address_inb = 123;
data_ina = 16'hffe6;
data_inb = 16'h6;
#10;
address_ina = 124;
address_inb = 125;
data_ina = 16'hfe74;
data_inb = 16'hfc1b;
#10;
address_ina = 126;
address_inb = 127;
data_ina = 16'h26f;
data_inb = 16'h333;
#10;
address_ina = 128;
address_inb = 129;
data_ina = 16'hffb9;
data_inb = 16'hfb71;
#10;
address_ina = 130;
address_inb = 131;
data_ina = 16'h47;
data_inb = 16'h535;
#10;
address_ina = 132;
address_inb = 133;
data_ina = 16'hfb15;
data_inb = 16'hfd76;
#10;
address_ina = 134;
address_inb = 135;
data_ina = 16'h13f;
data_inb = 16'h561;
#10;
address_ina = 136;
address_inb = 137;
data_ina = 16'hfef1;
data_inb = 16'hf990;
#10;
address_ina = 138;
address_inb = 139;
data_ina = 16'h67e;
data_inb = 16'hfb85;
#10;
address_ina = 140;
address_inb = 141;
data_ina = 16'hfa08;
data_inb = 16'hf9db;
#10;
address_ina = 142;
address_inb = 143;
data_ina = 16'hfda6;
data_inb = 16'h17b;
#10;
address_ina = 144;
address_inb = 145;
data_ina = 16'h103;
data_inb = 16'hf9fc;
#10;
address_ina = 146;
address_inb = 147;
data_ina = 16'hfacb;
data_inb = 16'hfcb1;
#10;
address_ina = 148;
address_inb = 149;
data_ina = 16'hfe9a;
data_inb = 16'hfeb7;
#10;
address_ina = 150;
address_inb = 151;
data_ina = 16'hffbc;
data_inb = 16'h397;
#10;
address_ina = 152;
address_inb = 153;
data_ina = 16'hf9fa;
data_inb = 16'h252;
#10;
address_ina = 154;
address_inb = 155;
data_ina = 16'hfd93;
data_inb = 16'hff32;
#10;
address_ina = 156;
address_inb = 157;
data_ina = 16'h596;
data_inb = 16'h478;
#10;
address_ina = 158;
address_inb = 159;
data_ina = 16'hfcaf;
data_inb = 16'h3e4;
#10;
address_ina = 160;
address_inb = 161;
data_ina = 16'h46a;
data_inb = 16'hfdde;
#10;
address_ina = 162;
address_inb = 163;
data_ina = 16'hf9a2;
data_inb = 16'h4de;
#10;
address_ina = 164;
address_inb = 165;
data_ina = 16'hfaf5;
data_inb = 16'h586;
#10;
address_ina = 166;
address_inb = 167;
data_ina = 16'hffbc;
data_inb = 16'hfc36;
#10;
address_ina = 168;
address_inb = 169;
data_ina = 16'hffd4;
data_inb = 16'h512;
#10;
address_ina = 170;
address_inb = 171;
data_ina = 16'hf9c9;
data_inb = 16'h19b;
#10;
address_ina = 172;
address_inb = 173;
data_ina = 16'h3e0;
data_inb = 16'hfccc;
#10;
address_ina = 174;
address_inb = 175;
data_ina = 16'h178;
data_inb = 16'h500;
#10;
address_ina = 176;
address_inb = 177;
data_ina = 16'hfb12;
data_inb = 16'hfd8c;
#10;
address_ina = 178;
address_inb = 179;
data_ina = 16'h3d5;
data_inb = 16'hfdff;
#10;
address_ina = 180;
address_inb = 181;
data_ina = 16'hfe66;
data_inb = 16'h42c;
#10;
address_ina = 182;
address_inb = 183;
data_ina = 16'hfa13;
data_inb = 16'hfa35;
#10;
address_ina = 184;
address_inb = 185;
data_ina = 16'hfc0d;
data_inb = 16'hfe91;
#10;
address_ina = 186;
address_inb = 187;
data_ina = 16'h5b7;
data_inb = 16'h357;
#10;
address_ina = 188;
address_inb = 189;
data_ina = 16'hbb;
data_inb = 16'hfcfb;
#10;
address_ina = 190;
address_inb = 191;
data_ina = 16'hfa7b;
data_inb = 16'h1ba;
#10;
address_ina = 192;
address_inb = 193;
data_ina = 16'hfada;
data_inb = 16'hfbf8;
#10;
address_ina = 194;
address_inb = 195;
data_ina = 16'h3ee;
data_inb = 16'h5d;
#10;
address_ina = 196;
address_inb = 197;
data_ina = 16'hf9da;
data_inb = 16'hfd4d;
#10;
address_ina = 198;
address_inb = 199;
data_ina = 16'hfbf5;
data_inb = 16'h11d;
#10;
address_ina = 200;
address_inb = 201;
data_ina = 16'hf988;
data_inb = 16'h4c0;
#10;
address_ina = 202;
address_inb = 203;
data_ina = 16'hfc38;
data_inb = 16'hfffa;
#10;
address_ina = 204;
address_inb = 205;
data_ina = 16'h262;
data_inb = 16'h5e6;
#10;
address_ina = 206;
address_inb = 207;
data_ina = 16'h137;
data_inb = 16'h307;
#10;
address_ina = 208;
address_inb = 209;
data_ina = 16'hfd3a;
data_inb = 16'h4b3;
#10;
address_ina = 210;
address_inb = 211;
data_ina = 16'hfd96;
data_inb = 16'hfccc;
#10;
address_ina = 212;
address_inb = 213;
data_ina = 16'hfc19;
data_inb = 16'hfce8;
#10;
address_ina = 214;
address_inb = 215;
data_ina = 16'h621;
data_inb = 16'h54b;
#10;
address_ina = 216;
address_inb = 217;
data_ina = 16'hfbc5;
data_inb = 16'h49e;
#10;
address_ina = 218;
address_inb = 219;
data_ina = 16'hfc1c;
data_inb = 16'hfd20;
#10;
address_ina = 220;
address_inb = 221;
data_ina = 16'h48f;
data_inb = 16'hfb62;
#10;
address_ina = 222;
address_inb = 223;
data_ina = 16'hfb61;
data_inb = 16'h570;
#10;
address_ina = 224;
address_inb = 225;
data_ina = 16'hfff5;
data_inb = 16'hfef5;
#10;
address_ina = 226;
address_inb = 227;
data_ina = 16'h380;
data_inb = 16'hf9ed;
#10;
address_ina = 228;
address_inb = 229;
data_ina = 16'h2d5;
data_inb = 16'h18a;
#10;
address_ina = 230;
address_inb = 231;
data_ina = 16'h2f1;
data_inb = 16'h657;
#10;
address_ina = 232;
address_inb = 233;
data_ina = 16'h4de;
data_inb = 16'hfd7a;
#10;
address_ina = 234;
address_inb = 235;
data_ina = 16'hfcad;
data_inb = 16'h37d;
#10;
address_ina = 236;
address_inb = 237;
data_ina = 16'h1e4;
data_inb = 16'h3d0;
#10;
address_ina = 238;
address_inb = 239;
data_ina = 16'h2b0;
data_inb = 16'hff54;
#10;
address_ina = 240;
address_inb = 241;
data_ina = 16'h34;
data_inb = 16'h504;
#10;
address_ina = 242;
address_inb = 243;
data_ina = 16'hfe8a;
data_inb = 16'h113;
#10;
address_ina = 244;
address_inb = 245;
data_ina = 16'hfde5;
data_inb = 16'hfa8d;
#10;
address_ina = 246;
address_inb = 247;
data_ina = 16'hfff7;
data_inb = 16'hff4f;
#10;
address_ina = 248;
address_inb = 249;
data_ina = 16'hffc4;
data_inb = 16'h409;
#10;
address_ina = 250;
address_inb = 251;
data_ina = 16'hf9cc;
data_inb = 16'hfd8b;
#10;
address_ina = 252;
address_inb = 253;
data_ina = 16'hfaec;
data_inb = 16'h5db;
#10;
address_ina = 254;
address_inb = 255;
data_ina = 16'hfed8;
data_inb = 16'h2a8;
#10;
        wait(init_done);
        #30
        we = 0;
        // Start processing
         
		  #38000

        start = 0;



//        wait (wr_req);
//		  wait (!wr_req);
//		   rd_req = 1;
		  wait(done);
		  #20000
rd_req = 1;
        #70 
		  start = 1;
		 #80 
wait(rd_empty)
rd_req = 0;

$display("Finished the NTT test Number %d",test_num);
////Begin test number #29//////////////
rst = 1;

//#1000
start = 1;
mode = 0; //NTT 0 // INTT 1

// Reset for a few clock cycles

#1000

rst = 0;
test_num = test_num + 1;
#1000
we = 1;
address_ina = 0;
address_inb = 1;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 2;
address_inb = 3;
data_ina = 16'h1;
data_inb = 16'h2;
#10;
address_ina = 4;
address_inb = 5;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 6;
address_inb = 7;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 8;
address_inb = 9;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 10;
address_inb = 11;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 12;
address_inb = 13;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 14;
address_inb = 15;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 16;
address_inb = 17;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 18;
address_inb = 19;
data_ina = 16'hfffe;
data_inb = 16'h1;
#10;
address_ina = 20;
address_inb = 21;
data_ina = 16'hfffe;
data_inb = 16'h1;
#10;
address_ina = 22;
address_inb = 23;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 24;
address_inb = 25;
data_ina = 16'h2;
data_inb = 16'h0;
#10;
address_ina = 26;
address_inb = 27;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 28;
address_inb = 29;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 30;
address_inb = 31;
data_ina = 16'hfffe;
data_inb = 16'h0;
#10;
address_ina = 32;
address_inb = 33;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 34;
address_inb = 35;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 36;
address_inb = 37;
data_ina = 16'hfffe;
data_inb = 16'hffff;
#10;
address_ina = 38;
address_inb = 39;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 40;
address_inb = 41;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 42;
address_inb = 43;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 44;
address_inb = 45;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 46;
address_inb = 47;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 48;
address_inb = 49;
data_ina = 16'hfffe;
data_inb = 16'h1;
#10;
address_ina = 50;
address_inb = 51;
data_ina = 16'h2;
data_inb = 16'hffff;
#10;
address_ina = 52;
address_inb = 53;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 54;
address_inb = 55;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 56;
address_inb = 57;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 58;
address_inb = 59;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 60;
address_inb = 61;
data_ina = 16'h0;
data_inb = 16'h2;
#10;
address_ina = 62;
address_inb = 63;
data_ina = 16'hfffe;
data_inb = 16'hffff;
#10;
address_ina = 64;
address_inb = 65;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 66;
address_inb = 67;
data_ina = 16'h3;
data_inb = 16'h0;
#10;
address_ina = 68;
address_inb = 69;
data_ina = 16'hffff;
data_inb = 16'hfffe;
#10;
address_ina = 70;
address_inb = 71;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 72;
address_inb = 73;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 74;
address_inb = 75;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 76;
address_inb = 77;
data_ina = 16'h2;
data_inb = 16'h2;
#10;
address_ina = 78;
address_inb = 79;
data_ina = 16'h2;
data_inb = 16'h0;
#10;
address_ina = 80;
address_inb = 81;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 82;
address_inb = 83;
data_ina = 16'h2;
data_inb = 16'h1;
#10;
address_ina = 84;
address_inb = 85;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 86;
address_inb = 87;
data_ina = 16'h0;
data_inb = 16'hfffe;
#10;
address_ina = 88;
address_inb = 89;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 90;
address_inb = 91;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 92;
address_inb = 93;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 94;
address_inb = 95;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 96;
address_inb = 97;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 98;
address_inb = 99;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 100;
address_inb = 101;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 102;
address_inb = 103;
data_ina = 16'h2;
data_inb = 16'h2;
#10;
address_ina = 104;
address_inb = 105;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 106;
address_inb = 107;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 108;
address_inb = 109;
data_ina = 16'h0;
data_inb = 16'h2;
#10;
address_ina = 110;
address_inb = 111;
data_ina = 16'h0;
data_inb = 16'hfffe;
#10;
address_ina = 112;
address_inb = 113;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 114;
address_inb = 115;
data_ina = 16'h0;
data_inb = 16'h2;
#10;
address_ina = 116;
address_inb = 117;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 118;
address_inb = 119;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 120;
address_inb = 121;
data_ina = 16'hffff;
data_inb = 16'hfffe;
#10;
address_ina = 122;
address_inb = 123;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 124;
address_inb = 125;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 126;
address_inb = 127;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 128;
address_inb = 129;
data_ina = 16'hfffd;
data_inb = 16'hffff;
#10;
address_ina = 130;
address_inb = 131;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 132;
address_inb = 133;
data_ina = 16'h0;
data_inb = 16'hfffd;
#10;
address_ina = 134;
address_inb = 135;
data_ina = 16'h0;
data_inb = 16'hfffe;
#10;
address_ina = 136;
address_inb = 137;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 138;
address_inb = 139;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 140;
address_inb = 141;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 142;
address_inb = 143;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 144;
address_inb = 145;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 146;
address_inb = 147;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 148;
address_inb = 149;
data_ina = 16'h1;
data_inb = 16'hfffe;
#10;
address_ina = 150;
address_inb = 151;
data_ina = 16'hffff;
data_inb = 16'h2;
#10;
address_ina = 152;
address_inb = 153;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 154;
address_inb = 155;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 156;
address_inb = 157;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 158;
address_inb = 159;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 160;
address_inb = 161;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 162;
address_inb = 163;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 164;
address_inb = 165;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 166;
address_inb = 167;
data_ina = 16'h0;
data_inb = 16'h2;
#10;
address_ina = 168;
address_inb = 169;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 170;
address_inb = 171;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 172;
address_inb = 173;
data_ina = 16'h0;
data_inb = 16'h2;
#10;
address_ina = 174;
address_inb = 175;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 176;
address_inb = 177;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 178;
address_inb = 179;
data_ina = 16'hfffe;
data_inb = 16'h1;
#10;
address_ina = 180;
address_inb = 181;
data_ina = 16'h2;
data_inb = 16'h2;
#10;
address_ina = 182;
address_inb = 183;
data_ina = 16'hfffe;
data_inb = 16'hffff;
#10;
address_ina = 184;
address_inb = 185;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 186;
address_inb = 187;
data_ina = 16'h3;
data_inb = 16'hffff;
#10;
address_ina = 188;
address_inb = 189;
data_ina = 16'h1;
data_inb = 16'h2;
#10;
address_ina = 190;
address_inb = 191;
data_ina = 16'h0;
data_inb = 16'hfffd;
#10;
address_ina = 192;
address_inb = 193;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 194;
address_inb = 195;
data_ina = 16'h2;
data_inb = 16'h0;
#10;
address_ina = 196;
address_inb = 197;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 198;
address_inb = 199;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 200;
address_inb = 201;
data_ina = 16'hfffe;
data_inb = 16'h1;
#10;
address_ina = 202;
address_inb = 203;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 204;
address_inb = 205;
data_ina = 16'h2;
data_inb = 16'h2;
#10;
address_ina = 206;
address_inb = 207;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 208;
address_inb = 209;
data_ina = 16'hfffe;
data_inb = 16'h2;
#10;
address_ina = 210;
address_inb = 211;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 212;
address_inb = 213;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 214;
address_inb = 215;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 216;
address_inb = 217;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 218;
address_inb = 219;
data_ina = 16'hfffe;
data_inb = 16'hfffe;
#10;
address_ina = 220;
address_inb = 221;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 222;
address_inb = 223;
data_ina = 16'h1;
data_inb = 16'hfffd;
#10;
address_ina = 224;
address_inb = 225;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 226;
address_inb = 227;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 228;
address_inb = 229;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 230;
address_inb = 231;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 232;
address_inb = 233;
data_ina = 16'h2;
data_inb = 16'h1;
#10;
address_ina = 234;
address_inb = 235;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 236;
address_inb = 237;
data_ina = 16'h0;
data_inb = 16'h2;
#10;
address_ina = 238;
address_inb = 239;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 240;
address_inb = 241;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 242;
address_inb = 243;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 244;
address_inb = 245;
data_ina = 16'h1;
data_inb = 16'h3;
#10;
address_ina = 246;
address_inb = 247;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 248;
address_inb = 249;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 250;
address_inb = 251;
data_ina = 16'hfffe;
data_inb = 16'h1;
#10;
address_ina = 252;
address_inb = 253;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 254;
address_inb = 255;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
        wait(init_done);
        #30
        we = 0;
        // Start processing
         
		  #38000

        start = 0;



//        wait (wr_req);
//		  wait (!wr_req);
//		   rd_req = 1;
		  wait(done);
		  #20000
rd_req = 1;
        #70 
		  start = 1;
		 #80 
wait(rd_empty)
rd_req = 0;

$display("Finished the NTT test Number %d",test_num);
////Begin test number #30//////////////
rst = 1;

//#1000
start = 1;
mode = 0; //NTT 0 // INTT 1

// Reset for a few clock cycles

#1000

rst = 0;
test_num = test_num + 1;
#1000
we = 1;
address_ina = 0;
address_inb = 1;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 2;
address_inb = 3;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 4;
address_inb = 5;
data_ina = 16'hfffe;
data_inb = 16'h2;
#10;
address_ina = 6;
address_inb = 7;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 8;
address_inb = 9;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 10;
address_inb = 11;
data_ina = 16'h2;
data_inb = 16'h0;
#10;
address_ina = 12;
address_inb = 13;
data_ina = 16'h2;
data_inb = 16'hfffe;
#10;
address_ina = 14;
address_inb = 15;
data_ina = 16'hfffe;
data_inb = 16'h1;
#10;
address_ina = 16;
address_inb = 17;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 18;
address_inb = 19;
data_ina = 16'hfffe;
data_inb = 16'h0;
#10;
address_ina = 20;
address_inb = 21;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 22;
address_inb = 23;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 24;
address_inb = 25;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 26;
address_inb = 27;
data_ina = 16'h2;
data_inb = 16'hffff;
#10;
address_ina = 28;
address_inb = 29;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 30;
address_inb = 31;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 32;
address_inb = 33;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 34;
address_inb = 35;
data_ina = 16'h2;
data_inb = 16'h1;
#10;
address_ina = 36;
address_inb = 37;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 38;
address_inb = 39;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 40;
address_inb = 41;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 42;
address_inb = 43;
data_ina = 16'hfffe;
data_inb = 16'hffff;
#10;
address_ina = 44;
address_inb = 45;
data_ina = 16'h1;
data_inb = 16'hfffe;
#10;
address_ina = 46;
address_inb = 47;
data_ina = 16'h2;
data_inb = 16'h0;
#10;
address_ina = 48;
address_inb = 49;
data_ina = 16'h0;
data_inb = 16'hfffe;
#10;
address_ina = 50;
address_inb = 51;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 52;
address_inb = 53;
data_ina = 16'hfffd;
data_inb = 16'hffff;
#10;
address_ina = 54;
address_inb = 55;
data_ina = 16'h1;
data_inb = 16'h2;
#10;
address_ina = 56;
address_inb = 57;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 58;
address_inb = 59;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 60;
address_inb = 61;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 62;
address_inb = 63;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 64;
address_inb = 65;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 66;
address_inb = 67;
data_ina = 16'h0;
data_inb = 16'hfffe;
#10;
address_ina = 68;
address_inb = 69;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 70;
address_inb = 71;
data_ina = 16'hffff;
data_inb = 16'hfffe;
#10;
address_ina = 72;
address_inb = 73;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 74;
address_inb = 75;
data_ina = 16'h0;
data_inb = 16'hfffe;
#10;
address_ina = 76;
address_inb = 77;
data_ina = 16'h2;
data_inb = 16'h0;
#10;
address_ina = 78;
address_inb = 79;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 80;
address_inb = 81;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 82;
address_inb = 83;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 84;
address_inb = 85;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 86;
address_inb = 87;
data_ina = 16'hffff;
data_inb = 16'h2;
#10;
address_ina = 88;
address_inb = 89;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 90;
address_inb = 91;
data_ina = 16'h0;
data_inb = 16'h2;
#10;
address_ina = 92;
address_inb = 93;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 94;
address_inb = 95;
data_ina = 16'hffff;
data_inb = 16'hfffe;
#10;
address_ina = 96;
address_inb = 97;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 98;
address_inb = 99;
data_ina = 16'h3;
data_inb = 16'hffff;
#10;
address_ina = 100;
address_inb = 101;
data_ina = 16'h0;
data_inb = 16'hfffe;
#10;
address_ina = 102;
address_inb = 103;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 104;
address_inb = 105;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 106;
address_inb = 107;
data_ina = 16'h0;
data_inb = 16'hfffe;
#10;
address_ina = 108;
address_inb = 109;
data_ina = 16'hfffd;
data_inb = 16'hfffe;
#10;
address_ina = 110;
address_inb = 111;
data_ina = 16'hfffd;
data_inb = 16'hffff;
#10;
address_ina = 112;
address_inb = 113;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 114;
address_inb = 115;
data_ina = 16'h0;
data_inb = 16'h2;
#10;
address_ina = 116;
address_inb = 117;
data_ina = 16'hffff;
data_inb = 16'hfffe;
#10;
address_ina = 118;
address_inb = 119;
data_ina = 16'hfffe;
data_inb = 16'h2;
#10;
address_ina = 120;
address_inb = 121;
data_ina = 16'h2;
data_inb = 16'hffff;
#10;
address_ina = 122;
address_inb = 123;
data_ina = 16'hffff;
data_inb = 16'h2;
#10;
address_ina = 124;
address_inb = 125;
data_ina = 16'h0;
data_inb = 16'h2;
#10;
address_ina = 126;
address_inb = 127;
data_ina = 16'hffff;
data_inb = 16'hfffe;
#10;
address_ina = 128;
address_inb = 129;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 130;
address_inb = 131;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 132;
address_inb = 133;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 134;
address_inb = 135;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 136;
address_inb = 137;
data_ina = 16'hfffe;
data_inb = 16'h0;
#10;
address_ina = 138;
address_inb = 139;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 140;
address_inb = 141;
data_ina = 16'hffff;
data_inb = 16'h2;
#10;
address_ina = 142;
address_inb = 143;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 144;
address_inb = 145;
data_ina = 16'h0;
data_inb = 16'hfffd;
#10;
address_ina = 146;
address_inb = 147;
data_ina = 16'h3;
data_inb = 16'h1;
#10;
address_ina = 148;
address_inb = 149;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 150;
address_inb = 151;
data_ina = 16'h2;
data_inb = 16'h0;
#10;
address_ina = 152;
address_inb = 153;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 154;
address_inb = 155;
data_ina = 16'h0;
data_inb = 16'h2;
#10;
address_ina = 156;
address_inb = 157;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 158;
address_inb = 159;
data_ina = 16'h2;
data_inb = 16'h2;
#10;
address_ina = 160;
address_inb = 161;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 162;
address_inb = 163;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 164;
address_inb = 165;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 166;
address_inb = 167;
data_ina = 16'h2;
data_inb = 16'h0;
#10;
address_ina = 168;
address_inb = 169;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 170;
address_inb = 171;
data_ina = 16'hfffd;
data_inb = 16'h1;
#10;
address_ina = 172;
address_inb = 173;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 174;
address_inb = 175;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 176;
address_inb = 177;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 178;
address_inb = 179;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 180;
address_inb = 181;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 182;
address_inb = 183;
data_ina = 16'h0;
data_inb = 16'hfffe;
#10;
address_ina = 184;
address_inb = 185;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 186;
address_inb = 187;
data_ina = 16'hfffe;
data_inb = 16'hfffd;
#10;
address_ina = 188;
address_inb = 189;
data_ina = 16'hfffe;
data_inb = 16'hffff;
#10;
address_ina = 190;
address_inb = 191;
data_ina = 16'h3;
data_inb = 16'h0;
#10;
address_ina = 192;
address_inb = 193;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 194;
address_inb = 195;
data_ina = 16'h2;
data_inb = 16'h0;
#10;
address_ina = 196;
address_inb = 197;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 198;
address_inb = 199;
data_ina = 16'h2;
data_inb = 16'h2;
#10;
address_ina = 200;
address_inb = 201;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 202;
address_inb = 203;
data_ina = 16'hfffd;
data_inb = 16'hffff;
#10;
address_ina = 204;
address_inb = 205;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 206;
address_inb = 207;
data_ina = 16'hfffe;
data_inb = 16'hffff;
#10;
address_ina = 208;
address_inb = 209;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 210;
address_inb = 211;
data_ina = 16'h0;
data_inb = 16'hfffe;
#10;
address_ina = 212;
address_inb = 213;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 214;
address_inb = 215;
data_ina = 16'hfffe;
data_inb = 16'h0;
#10;
address_ina = 216;
address_inb = 217;
data_ina = 16'h1;
data_inb = 16'h2;
#10;
address_ina = 218;
address_inb = 219;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 220;
address_inb = 221;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 222;
address_inb = 223;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 224;
address_inb = 225;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 226;
address_inb = 227;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 228;
address_inb = 229;
data_ina = 16'hffff;
data_inb = 16'hfffe;
#10;
address_ina = 230;
address_inb = 231;
data_ina = 16'hfffe;
data_inb = 16'hfffe;
#10;
address_ina = 232;
address_inb = 233;
data_ina = 16'hffff;
data_inb = 16'h2;
#10;
address_ina = 234;
address_inb = 235;
data_ina = 16'hffff;
data_inb = 16'hfffe;
#10;
address_ina = 236;
address_inb = 237;
data_ina = 16'hffff;
data_inb = 16'h2;
#10;
address_ina = 238;
address_inb = 239;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 240;
address_inb = 241;
data_ina = 16'h3;
data_inb = 16'h1;
#10;
address_ina = 242;
address_inb = 243;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 244;
address_inb = 245;
data_ina = 16'hfffe;
data_inb = 16'h1;
#10;
address_ina = 246;
address_inb = 247;
data_ina = 16'hfffe;
data_inb = 16'hffff;
#10;
address_ina = 248;
address_inb = 249;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 250;
address_inb = 251;
data_ina = 16'hffff;
data_inb = 16'h2;
#10;
address_ina = 252;
address_inb = 253;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 254;
address_inb = 255;
data_ina = 16'h1;
data_inb = 16'hfffe;
#10;
        wait(init_done);
        #30
        we = 0;
        // Start processing
         
		  #38000

        start = 0;



//        wait (wr_req);
//		  wait (!wr_req);
//		   rd_req = 1;
		  wait(done);
		  #20000
rd_req = 1;
        #70 
		  start = 1;
		 #80 
wait(rd_empty)
rd_req = 0;

$display("Finished the NTT test Number %d",test_num);
////Begin test number #31//////////////
rst = 1;

//#1000
start = 1;
mode = 1; //NTT 0 // INTT 1

// Reset for a few clock cycles

#1000

rst = 0;
test_num = test_num + 1;
#1000
we = 1;
address_ina = 0;
address_inb = 1;
data_ina = 16'hfc65;
data_inb = 16'h88;
#10;
address_ina = 2;
address_inb = 3;
data_ina = 16'h5e7;
data_inb = 16'h30f;
#10;
address_ina = 4;
address_inb = 5;
data_ina = 16'h3f6;
data_inb = 16'h47f;
#10;
address_ina = 6;
address_inb = 7;
data_ina = 16'hfd0a;
data_inb = 16'h3c6;
#10;
address_ina = 8;
address_inb = 9;
data_ina = 16'hfc6c;
data_inb = 16'he5;
#10;
address_ina = 10;
address_inb = 11;
data_ina = 16'h29b;
data_inb = 16'hfd98;
#10;
address_ina = 12;
address_inb = 13;
data_ina = 16'hf9c2;
data_inb = 16'hfac6;
#10;
address_ina = 14;
address_inb = 15;
data_ina = 16'hfcfb;
data_inb = 16'h419;
#10;
address_ina = 16;
address_inb = 17;
data_ina = 16'hffd7;
data_inb = 16'h42f;
#10;
address_ina = 18;
address_inb = 19;
data_ina = 16'h24a;
data_inb = 16'h15f;
#10;
address_ina = 20;
address_inb = 21;
data_ina = 16'hfe1a;
data_inb = 16'h560;
#10;
address_ina = 22;
address_inb = 23;
data_ina = 16'hff82;
data_inb = 16'hfcf9;
#10;
address_ina = 24;
address_inb = 25;
data_ina = 16'h103;
data_inb = 16'hfac3;
#10;
address_ina = 26;
address_inb = 27;
data_ina = 16'h2f;
data_inb = 16'h2df;
#10;
address_ina = 28;
address_inb = 29;
data_ina = 16'h36d;
data_inb = 16'hfccc;
#10;
address_ina = 30;
address_inb = 31;
data_ina = 16'h197;
data_inb = 16'hfdcc;
#10;
address_ina = 32;
address_inb = 33;
data_ina = 16'hfa23;
data_inb = 16'h214;
#10;
address_ina = 34;
address_inb = 35;
data_ina = 16'h35;
data_inb = 16'hfdb2;
#10;
address_ina = 36;
address_inb = 37;
data_ina = 16'h47e;
data_inb = 16'h6b;
#10;
address_ina = 38;
address_inb = 39;
data_ina = 16'hfa0d;
data_inb = 16'h62;
#10;
address_ina = 40;
address_inb = 41;
data_ina = 16'h3b5;
data_inb = 16'h401;
#10;
address_ina = 42;
address_inb = 43;
data_ina = 16'hfe0b;
data_inb = 16'h5a2;
#10;
address_ina = 44;
address_inb = 45;
data_ina = 16'h95;
data_inb = 16'hfff6;
#10;
address_ina = 46;
address_inb = 47;
data_ina = 16'h143;
data_inb = 16'h2c9;
#10;
address_ina = 48;
address_inb = 49;
data_ina = 16'hfe04;
data_inb = 16'h23a;
#10;
address_ina = 50;
address_inb = 51;
data_ina = 16'h380;
data_inb = 16'h4e4;
#10;
address_ina = 52;
address_inb = 53;
data_ina = 16'h356;
data_inb = 16'h128;
#10;
address_ina = 54;
address_inb = 55;
data_ina = 16'h4c3;
data_inb = 16'h3c8;
#10;
address_ina = 56;
address_inb = 57;
data_ina = 16'h1ab;
data_inb = 16'h547;
#10;
address_ina = 58;
address_inb = 59;
data_ina = 16'hfa7c;
data_inb = 16'hfa9f;
#10;
address_ina = 60;
address_inb = 61;
data_ina = 16'hfe49;
data_inb = 16'h536;
#10;
address_ina = 62;
address_inb = 63;
data_ina = 16'h30e;
data_inb = 16'h51f;
#10;
address_ina = 64;
address_inb = 65;
data_ina = 16'hfd98;
data_inb = 16'hffff;
#10;
address_ina = 66;
address_inb = 67;
data_ina = 16'h36;
data_inb = 16'h5c7;
#10;
address_ina = 68;
address_inb = 69;
data_ina = 16'h1c4;
data_inb = 16'h1cb;
#10;
address_ina = 70;
address_inb = 71;
data_ina = 16'h454;
data_inb = 16'h415;
#10;
address_ina = 72;
address_inb = 73;
data_ina = 16'h5fa;
data_inb = 16'h596;
#10;
address_ina = 74;
address_inb = 75;
data_ina = 16'hfcd2;
data_inb = 16'hfb9c;
#10;
address_ina = 76;
address_inb = 77;
data_ina = 16'hffff;
data_inb = 16'h58f;
#10;
address_ina = 78;
address_inb = 79;
data_ina = 16'hfdae;
data_inb = 16'h60e;
#10;
address_ina = 80;
address_inb = 81;
data_ina = 16'h34a;
data_inb = 16'h29;
#10;
address_ina = 82;
address_inb = 83;
data_ina = 16'h650;
data_inb = 16'hfb15;
#10;
address_ina = 84;
address_inb = 85;
data_ina = 16'hfd7c;
data_inb = 16'hfc21;
#10;
address_ina = 86;
address_inb = 87;
data_ina = 16'h658;
data_inb = 16'h627;
#10;
address_ina = 88;
address_inb = 89;
data_ina = 16'h4c2;
data_inb = 16'hfe6d;
#10;
address_ina = 90;
address_inb = 91;
data_ina = 16'hff01;
data_inb = 16'hfb8d;
#10;
address_ina = 92;
address_inb = 93;
data_ina = 16'hfe9e;
data_inb = 16'hf9fc;
#10;
address_ina = 94;
address_inb = 95;
data_ina = 16'hf9ef;
data_inb = 16'hfb1d;
#10;
address_ina = 96;
address_inb = 97;
data_ina = 16'h43d;
data_inb = 16'hfc10;
#10;
address_ina = 98;
address_inb = 99;
data_ina = 16'h300;
data_inb = 16'h609;
#10;
address_ina = 100;
address_inb = 101;
data_ina = 16'hab;
data_inb = 16'hfbe1;
#10;
address_ina = 102;
address_inb = 103;
data_ina = 16'hfdd5;
data_inb = 16'hfd36;
#10;
address_ina = 104;
address_inb = 105;
data_ina = 16'h35e;
data_inb = 16'hfb0c;
#10;
address_ina = 106;
address_inb = 107;
data_ina = 16'h10a;
data_inb = 16'hfe25;
#10;
address_ina = 108;
address_inb = 109;
data_ina = 16'hfc6c;
data_inb = 16'hfbeb;
#10;
address_ina = 110;
address_inb = 111;
data_ina = 16'hfc6f;
data_inb = 16'h1b4;
#10;
address_ina = 112;
address_inb = 113;
data_ina = 16'hfaf0;
data_inb = 16'h2c7;
#10;
address_ina = 114;
address_inb = 115;
data_ina = 16'hfc50;
data_inb = 16'h2ec;
#10;
address_ina = 116;
address_inb = 117;
data_ina = 16'h46c;
data_inb = 16'h67f;
#10;
address_ina = 118;
address_inb = 119;
data_ina = 16'ha9;
data_inb = 16'h304;
#10;
address_ina = 120;
address_inb = 121;
data_ina = 16'hba;
data_inb = 16'h5b6;
#10;
address_ina = 122;
address_inb = 123;
data_ina = 16'hfe79;
data_inb = 16'h412;
#10;
address_ina = 124;
address_inb = 125;
data_ina = 16'hffcf;
data_inb = 16'h2cd;
#10;
address_ina = 126;
address_inb = 127;
data_ina = 16'hfc5b;
data_inb = 16'hfe45;
#10;
address_ina = 128;
address_inb = 129;
data_ina = 16'h3f8;
data_inb = 16'h357;
#10;
address_ina = 130;
address_inb = 131;
data_ina = 16'hff85;
data_inb = 16'hff57;
#10;
address_ina = 132;
address_inb = 133;
data_ina = 16'hfb76;
data_inb = 16'hf9c0;
#10;
address_ina = 134;
address_inb = 135;
data_ina = 16'hff70;
data_inb = 16'h11;
#10;
address_ina = 136;
address_inb = 137;
data_ina = 16'hfffe;
data_inb = 16'hfe20;
#10;
address_ina = 138;
address_inb = 139;
data_ina = 16'hfec5;
data_inb = 16'hfe31;
#10;
address_ina = 140;
address_inb = 141;
data_ina = 16'h3cd;
data_inb = 16'h352;
#10;
address_ina = 142;
address_inb = 143;
data_ina = 16'h5bc;
data_inb = 16'hfb33;
#10;
address_ina = 144;
address_inb = 145;
data_ina = 16'hfe6a;
data_inb = 16'hfc4d;
#10;
address_ina = 146;
address_inb = 147;
data_ina = 16'h418;
data_inb = 16'h5d2;
#10;
address_ina = 148;
address_inb = 149;
data_ina = 16'h36a;
data_inb = 16'hfe00;
#10;
address_ina = 150;
address_inb = 151;
data_ina = 16'h38d;
data_inb = 16'h2c8;
#10;
address_ina = 152;
address_inb = 153;
data_ina = 16'h2a4;
data_inb = 16'hfe68;
#10;
address_ina = 154;
address_inb = 155;
data_ina = 16'h37d;
data_inb = 16'h435;
#10;
address_ina = 156;
address_inb = 157;
data_ina = 16'h50c;
data_inb = 16'h632;
#10;
address_ina = 158;
address_inb = 159;
data_ina = 16'h43b;
data_inb = 16'h461;
#10;
address_ina = 160;
address_inb = 161;
data_ina = 16'hffb0;
data_inb = 16'hfa8b;
#10;
address_ina = 162;
address_inb = 163;
data_ina = 16'h211;
data_inb = 16'hffa3;
#10;
address_ina = 164;
address_inb = 165;
data_ina = 16'h507;
data_inb = 16'h4f5;
#10;
address_ina = 166;
address_inb = 167;
data_ina = 16'hfab8;
data_inb = 16'hfc84;
#10;
address_ina = 168;
address_inb = 169;
data_ina = 16'h198;
data_inb = 16'hfbdb;
#10;
address_ina = 170;
address_inb = 171;
data_ina = 16'h567;
data_inb = 16'hfe33;
#10;
address_ina = 172;
address_inb = 173;
data_ina = 16'hc1;
data_inb = 16'h58b;
#10;
address_ina = 174;
address_inb = 175;
data_ina = 16'hfc1f;
data_inb = 16'h58;
#10;
address_ina = 176;
address_inb = 177;
data_ina = 16'hfd9f;
data_inb = 16'hfeed;
#10;
address_ina = 178;
address_inb = 179;
data_ina = 16'h128;
data_inb = 16'hfdc9;
#10;
address_ina = 180;
address_inb = 181;
data_ina = 16'hfd41;
data_inb = 16'hfbc6;
#10;
address_ina = 182;
address_inb = 183;
data_ina = 16'h2c2;
data_inb = 16'h0;
#10;
address_ina = 184;
address_inb = 185;
data_ina = 16'hfb5f;
data_inb = 16'hfe7a;
#10;
address_ina = 186;
address_inb = 187;
data_ina = 16'hff6c;
data_inb = 16'hfd9b;
#10;
address_ina = 188;
address_inb = 189;
data_ina = 16'hfa2e;
data_inb = 16'h453;
#10;
address_ina = 190;
address_inb = 191;
data_ina = 16'h2e1;
data_inb = 16'h5b4;
#10;
address_ina = 192;
address_inb = 193;
data_ina = 16'hffed;
data_inb = 16'hfe0e;
#10;
address_ina = 194;
address_inb = 195;
data_ina = 16'h35a;
data_inb = 16'h2ff;
#10;
address_ina = 196;
address_inb = 197;
data_ina = 16'hff26;
data_inb = 16'hff28;
#10;
address_ina = 198;
address_inb = 199;
data_ina = 16'hfcff;
data_inb = 16'haa;
#10;
address_ina = 200;
address_inb = 201;
data_ina = 16'h1f;
data_inb = 16'h228;
#10;
address_ina = 202;
address_inb = 203;
data_ina = 16'hfe1c;
data_inb = 16'hfbe3;
#10;
address_ina = 204;
address_inb = 205;
data_ina = 16'h1b2;
data_inb = 16'h63a;
#10;
address_ina = 206;
address_inb = 207;
data_ina = 16'h560;
data_inb = 16'hfc46;
#10;
address_ina = 208;
address_inb = 209;
data_ina = 16'h257;
data_inb = 16'h150;
#10;
address_ina = 210;
address_inb = 211;
data_ina = 16'hfe65;
data_inb = 16'h231;
#10;
address_ina = 212;
address_inb = 213;
data_ina = 16'hf9b2;
data_inb = 16'hfa10;
#10;
address_ina = 214;
address_inb = 215;
data_ina = 16'h499;
data_inb = 16'hfa39;
#10;
address_ina = 216;
address_inb = 217;
data_ina = 16'hfd87;
data_inb = 16'h2ef;
#10;
address_ina = 218;
address_inb = 219;
data_ina = 16'hc7;
data_inb = 16'h190;
#10;
address_ina = 220;
address_inb = 221;
data_ina = 16'h5ab;
data_inb = 16'hfa4c;
#10;
address_ina = 222;
address_inb = 223;
data_ina = 16'hfd;
data_inb = 16'h420;
#10;
address_ina = 224;
address_inb = 225;
data_ina = 16'h284;
data_inb = 16'hffe0;
#10;
address_ina = 226;
address_inb = 227;
data_ina = 16'h2a2;
data_inb = 16'h437;
#10;
address_ina = 228;
address_inb = 229;
data_ina = 16'h413;
data_inb = 16'hfda8;
#10;
address_ina = 230;
address_inb = 231;
data_ina = 16'hfe2c;
data_inb = 16'h11;
#10;
address_ina = 232;
address_inb = 233;
data_ina = 16'hf9d0;
data_inb = 16'hfcbe;
#10;
address_ina = 234;
address_inb = 235;
data_ina = 16'h464;
data_inb = 16'h1e4;
#10;
address_ina = 236;
address_inb = 237;
data_ina = 16'h2b;
data_inb = 16'hfce8;
#10;
address_ina = 238;
address_inb = 239;
data_ina = 16'hfda4;
data_inb = 16'hff2d;
#10;
address_ina = 240;
address_inb = 241;
data_ina = 16'hfa5a;
data_inb = 16'h9d;
#10;
address_ina = 242;
address_inb = 243;
data_ina = 16'h5c1;
data_inb = 16'hfe21;
#10;
address_ina = 244;
address_inb = 245;
data_ina = 16'hfd8e;
data_inb = 16'hfc83;
#10;
address_ina = 246;
address_inb = 247;
data_ina = 16'hff65;
data_inb = 16'h341;
#10;
address_ina = 248;
address_inb = 249;
data_ina = 16'h7f;
data_inb = 16'hfb4d;
#10;
address_ina = 250;
address_inb = 251;
data_ina = 16'h332;
data_inb = 16'h528;
#10;
address_ina = 252;
address_inb = 253;
data_ina = 16'hfdec;
data_inb = 16'hfbe6;
#10;
address_ina = 254;
address_inb = 255;
data_ina = 16'hfed0;
data_inb = 16'hfd3e;
#10;
        wait(init_done);
        #30
        we = 0;
        // Start processing
         
		  #38000

        start = 0;



//        wait (wr_req);
//		  wait (!wr_req);
//		   rd_req = 1;
		  wait(done);
		  #20000
rd_req = 1;
        #70 
		  start = 1;
		 #80 
wait(rd_empty)
rd_req = 0;

$display("Finished the NTT test Number %d",test_num);
////Begin test number #32//////////////
rst = 1;

//#1000
start = 1;
mode = 1; //NTT 0 // INTT 1

// Reset for a few clock cycles

#1000

rst = 0;
test_num = test_num + 1;
#1000
we = 1;
address_ina = 0;
address_inb = 1;
data_ina = 16'h13c;
data_inb = 16'hfd50;
#10;
address_ina = 2;
address_inb = 3;
data_ina = 16'hf9e0;
data_inb = 16'hfba0;
#10;
address_ina = 4;
address_inb = 5;
data_ina = 16'h629;
data_inb = 16'h541;
#10;
address_ina = 6;
address_inb = 7;
data_ina = 16'h608;
data_inb = 16'hff9c;
#10;
address_ina = 8;
address_inb = 9;
data_ina = 16'h149;
data_inb = 16'h288;
#10;
address_ina = 10;
address_inb = 11;
data_ina = 16'hfcdd;
data_inb = 16'h249;
#10;
address_ina = 12;
address_inb = 13;
data_ina = 16'hfc44;
data_inb = 16'hfaf7;
#10;
address_ina = 14;
address_inb = 15;
data_ina = 16'h172;
data_inb = 16'h359;
#10;
address_ina = 16;
address_inb = 17;
data_ina = 16'h35d;
data_inb = 16'hfb0b;
#10;
address_ina = 18;
address_inb = 19;
data_ina = 16'hfdec;
data_inb = 16'h115;
#10;
address_ina = 20;
address_inb = 21;
data_ina = 16'h424;
data_inb = 16'hfffd;
#10;
address_ina = 22;
address_inb = 23;
data_ina = 16'hfe1f;
data_inb = 16'hfb56;
#10;
address_ina = 24;
address_inb = 25;
data_ina = 16'hfa4f;
data_inb = 16'hfca0;
#10;
address_ina = 26;
address_inb = 27;
data_ina = 16'h3df;
data_inb = 16'hffc8;
#10;
address_ina = 28;
address_inb = 29;
data_ina = 16'h4ed;
data_inb = 16'hfdff;
#10;
address_ina = 30;
address_inb = 31;
data_ina = 16'hfdf6;
data_inb = 16'hfd18;
#10;
address_ina = 32;
address_inb = 33;
data_ina = 16'hfd0a;
data_inb = 16'h477;
#10;
address_ina = 34;
address_inb = 35;
data_ina = 16'h19a;
data_inb = 16'hfdf0;
#10;
address_ina = 36;
address_inb = 37;
data_ina = 16'hfa22;
data_inb = 16'h26c;
#10;
address_ina = 38;
address_inb = 39;
data_ina = 16'hfe5d;
data_inb = 16'hfca9;
#10;
address_ina = 40;
address_inb = 41;
data_ina = 16'h9d;
data_inb = 16'hffe1;
#10;
address_ina = 42;
address_inb = 43;
data_ina = 16'hfbff;
data_inb = 16'h196;
#10;
address_ina = 44;
address_inb = 45;
data_ina = 16'h3ac;
data_inb = 16'hfd4c;
#10;
address_ina = 46;
address_inb = 47;
data_ina = 16'h1c3;
data_inb = 16'hfe60;
#10;
address_ina = 48;
address_inb = 49;
data_ina = 16'hfa55;
data_inb = 16'h30b;
#10;
address_ina = 50;
address_inb = 51;
data_ina = 16'hff30;
data_inb = 16'hfbbc;
#10;
address_ina = 52;
address_inb = 53;
data_ina = 16'hff90;
data_inb = 16'h287;
#10;
address_ina = 54;
address_inb = 55;
data_ina = 16'h5ec;
data_inb = 16'hf99e;
#10;
address_ina = 56;
address_inb = 57;
data_ina = 16'hba;
data_inb = 16'hfc15;
#10;
address_ina = 58;
address_inb = 59;
data_ina = 16'h2f7;
data_inb = 16'hbb;
#10;
address_ina = 60;
address_inb = 61;
data_ina = 16'hfcd8;
data_inb = 16'h37e;
#10;
address_ina = 62;
address_inb = 63;
data_ina = 16'hf9ce;
data_inb = 16'h4b4;
#10;
address_ina = 64;
address_inb = 65;
data_ina = 16'h615;
data_inb = 16'h472;
#10;
address_ina = 66;
address_inb = 67;
data_ina = 16'hf997;
data_inb = 16'hfd85;
#10;
address_ina = 68;
address_inb = 69;
data_ina = 16'h295;
data_inb = 16'hfaf8;
#10;
address_ina = 70;
address_inb = 71;
data_ina = 16'h136;
data_inb = 16'hf986;
#10;
address_ina = 72;
address_inb = 73;
data_ina = 16'h1c6;
data_inb = 16'h477;
#10;
address_ina = 74;
address_inb = 75;
data_ina = 16'h1fe;
data_inb = 16'hfa2c;
#10;
address_ina = 76;
address_inb = 77;
data_ina = 16'hfceb;
data_inb = 16'h443;
#10;
address_ina = 78;
address_inb = 79;
data_ina = 16'h66c;
data_inb = 16'hffc3;
#10;
address_ina = 80;
address_inb = 81;
data_ina = 16'hfdc0;
data_inb = 16'hfb1a;
#10;
address_ina = 82;
address_inb = 83;
data_ina = 16'h11;
data_inb = 16'h119;
#10;
address_ina = 84;
address_inb = 85;
data_ina = 16'hfc57;
data_inb = 16'h644;
#10;
address_ina = 86;
address_inb = 87;
data_ina = 16'h13b;
data_inb = 16'h51a;
#10;
address_ina = 88;
address_inb = 89;
data_ina = 16'hfc65;
data_inb = 16'hfa5b;
#10;
address_ina = 90;
address_inb = 91;
data_ina = 16'h4fd;
data_inb = 16'hf982;
#10;
address_ina = 92;
address_inb = 93;
data_ina = 16'h374;
data_inb = 16'h59b;
#10;
address_ina = 94;
address_inb = 95;
data_ina = 16'hfa3b;
data_inb = 16'h3c2;
#10;
address_ina = 96;
address_inb = 97;
data_ina = 16'hfc73;
data_inb = 16'h20c;
#10;
address_ina = 98;
address_inb = 99;
data_ina = 16'h296;
data_inb = 16'hfb5f;
#10;
address_ina = 100;
address_inb = 101;
data_ina = 16'h557;
data_inb = 16'h2a5;
#10;
address_ina = 102;
address_inb = 103;
data_ina = 16'hfded;
data_inb = 16'h3b5;
#10;
address_ina = 104;
address_inb = 105;
data_ina = 16'hfd2b;
data_inb = 16'h4cb;
#10;
address_ina = 106;
address_inb = 107;
data_ina = 16'h4f2;
data_inb = 16'h634;
#10;
address_ina = 108;
address_inb = 109;
data_ina = 16'h573;
data_inb = 16'h18f;
#10;
address_ina = 110;
address_inb = 111;
data_ina = 16'h60f;
data_inb = 16'h1fa;
#10;
address_ina = 112;
address_inb = 113;
data_ina = 16'h1c6;
data_inb = 16'hfcc4;
#10;
address_ina = 114;
address_inb = 115;
data_ina = 16'hfcd1;
data_inb = 16'h55f;
#10;
address_ina = 116;
address_inb = 117;
data_ina = 16'h390;
data_inb = 16'h22a;
#10;
address_ina = 118;
address_inb = 119;
data_ina = 16'h36f;
data_inb = 16'hfe21;
#10;
address_ina = 120;
address_inb = 121;
data_ina = 16'h370;
data_inb = 16'h126;
#10;
address_ina = 122;
address_inb = 123;
data_ina = 16'hfb44;
data_inb = 16'hfa8d;
#10;
address_ina = 124;
address_inb = 125;
data_ina = 16'h17d;
data_inb = 16'hfe7c;
#10;
address_ina = 126;
address_inb = 127;
data_ina = 16'h4e7;
data_inb = 16'hfe84;
#10;
address_ina = 128;
address_inb = 129;
data_ina = 16'hfa8e;
data_inb = 16'hfe3b;
#10;
address_ina = 130;
address_inb = 131;
data_ina = 16'hfe03;
data_inb = 16'h3b5;
#10;
address_ina = 132;
address_inb = 133;
data_ina = 16'h3ed;
data_inb = 16'h37f;
#10;
address_ina = 134;
address_inb = 135;
data_ina = 16'hff0b;
data_inb = 16'ha7;
#10;
address_ina = 136;
address_inb = 137;
data_ina = 16'h17d;
data_inb = 16'h18d;
#10;
address_ina = 138;
address_inb = 139;
data_ina = 16'hffcf;
data_inb = 16'h5ba;
#10;
address_ina = 140;
address_inb = 141;
data_ina = 16'hfea2;
data_inb = 16'h457;
#10;
address_ina = 142;
address_inb = 143;
data_ina = 16'h13d;
data_inb = 16'h10d;
#10;
address_ina = 144;
address_inb = 145;
data_ina = 16'h5cc;
data_inb = 16'h2ef;
#10;
address_ina = 146;
address_inb = 147;
data_ina = 16'hfec6;
data_inb = 16'h19c;
#10;
address_ina = 148;
address_inb = 149;
data_ina = 16'hfaf4;
data_inb = 16'hfb84;
#10;
address_ina = 150;
address_inb = 151;
data_ina = 16'h131;
data_inb = 16'h475;
#10;
address_ina = 152;
address_inb = 153;
data_ina = 16'h116;
data_inb = 16'hfa79;
#10;
address_ina = 154;
address_inb = 155;
data_ina = 16'h3b2;
data_inb = 16'hff9b;
#10;
address_ina = 156;
address_inb = 157;
data_ina = 16'hfafb;
data_inb = 16'h37b;
#10;
address_ina = 158;
address_inb = 159;
data_ina = 16'hfb33;
data_inb = 16'hfd76;
#10;
address_ina = 160;
address_inb = 161;
data_ina = 16'h198;
data_inb = 16'h478;
#10;
address_ina = 162;
address_inb = 163;
data_ina = 16'h66d;
data_inb = 16'h406;
#10;
address_ina = 164;
address_inb = 165;
data_ina = 16'h5ca;
data_inb = 16'hffe6;
#10;
address_ina = 166;
address_inb = 167;
data_ina = 16'h61;
data_inb = 16'h3;
#10;
address_ina = 168;
address_inb = 169;
data_ina = 16'h1df;
data_inb = 16'hfff0;
#10;
address_ina = 170;
address_inb = 171;
data_ina = 16'hfb63;
data_inb = 16'hfffb;
#10;
address_ina = 172;
address_inb = 173;
data_ina = 16'h1d2;
data_inb = 16'hfc6e;
#10;
address_ina = 174;
address_inb = 175;
data_ina = 16'h27b;
data_inb = 16'hfd5b;
#10;
address_ina = 176;
address_inb = 177;
data_ina = 16'hfc1e;
data_inb = 16'hfe0f;
#10;
address_ina = 178;
address_inb = 179;
data_ina = 16'h27b;
data_inb = 16'hfd45;
#10;
address_ina = 180;
address_inb = 181;
data_ina = 16'hfdef;
data_inb = 16'h21c;
#10;
address_ina = 182;
address_inb = 183;
data_ina = 16'h5af;
data_inb = 16'hfb75;
#10;
address_ina = 184;
address_inb = 185;
data_ina = 16'hfaec;
data_inb = 16'hfd6d;
#10;
address_ina = 186;
address_inb = 187;
data_ina = 16'h106;
data_inb = 16'hfe91;
#10;
address_ina = 188;
address_inb = 189;
data_ina = 16'h4f4;
data_inb = 16'h3f1;
#10;
address_ina = 190;
address_inb = 191;
data_ina = 16'h5a1;
data_inb = 16'h1da;
#10;
address_ina = 192;
address_inb = 193;
data_ina = 16'h2ee;
data_inb = 16'hfde8;
#10;
address_ina = 194;
address_inb = 195;
data_ina = 16'h1a3;
data_inb = 16'hfe52;
#10;
address_ina = 196;
address_inb = 197;
data_ina = 16'hfd47;
data_inb = 16'hfd19;
#10;
address_ina = 198;
address_inb = 199;
data_ina = 16'hffbc;
data_inb = 16'hfbc3;
#10;
address_ina = 200;
address_inb = 201;
data_ina = 16'h1ef;
data_inb = 16'hfd80;
#10;
address_ina = 202;
address_inb = 203;
data_ina = 16'h222;
data_inb = 16'hd;
#10;
address_ina = 204;
address_inb = 205;
data_ina = 16'hff66;
data_inb = 16'hfd55;
#10;
address_ina = 206;
address_inb = 207;
data_ina = 16'hfbc8;
data_inb = 16'hfccc;
#10;
address_ina = 208;
address_inb = 209;
data_ina = 16'h4d0;
data_inb = 16'h43e;
#10;
address_ina = 210;
address_inb = 211;
data_ina = 16'h49f;
data_inb = 16'hfdcf;
#10;
address_ina = 212;
address_inb = 213;
data_ina = 16'h2fb;
data_inb = 16'h5cd;
#10;
address_ina = 214;
address_inb = 215;
data_ina = 16'hfb5f;
data_inb = 16'hfbec;
#10;
address_ina = 216;
address_inb = 217;
data_ina = 16'hfe74;
data_inb = 16'h374;
#10;
address_ina = 218;
address_inb = 219;
data_ina = 16'hff21;
data_inb = 16'hf5;
#10;
address_ina = 220;
address_inb = 221;
data_ina = 16'hfad9;
data_inb = 16'hfe06;
#10;
address_ina = 222;
address_inb = 223;
data_ina = 16'h1b1;
data_inb = 16'h55e;
#10;
address_ina = 224;
address_inb = 225;
data_ina = 16'h109;
data_inb = 16'hfd85;
#10;
address_ina = 226;
address_inb = 227;
data_ina = 16'h604;
data_inb = 16'hfb3d;
#10;
address_ina = 228;
address_inb = 229;
data_ina = 16'hf987;
data_inb = 16'hfb8c;
#10;
address_ina = 230;
address_inb = 231;
data_ina = 16'h4e0;
data_inb = 16'hf9b5;
#10;
address_ina = 232;
address_inb = 233;
data_ina = 16'hfc53;
data_inb = 16'hfaed;
#10;
address_ina = 234;
address_inb = 235;
data_ina = 16'h1f3;
data_inb = 16'hfe50;
#10;
address_ina = 236;
address_inb = 237;
data_ina = 16'hfcf5;
data_inb = 16'h52f;
#10;
address_ina = 238;
address_inb = 239;
data_ina = 16'hff43;
data_inb = 16'h1fc;
#10;
address_ina = 240;
address_inb = 241;
data_ina = 16'h15e;
data_inb = 16'h1b1;
#10;
address_ina = 242;
address_inb = 243;
data_ina = 16'h343;
data_inb = 16'hfa8a;
#10;
address_ina = 244;
address_inb = 245;
data_ina = 16'hfbaa;
data_inb = 16'h53c;
#10;
address_ina = 246;
address_inb = 247;
data_ina = 16'h26b;
data_inb = 16'hfd0c;
#10;
address_ina = 248;
address_inb = 249;
data_ina = 16'h15f;
data_inb = 16'hfe6a;
#10;
address_ina = 250;
address_inb = 251;
data_ina = 16'hf0;
data_inb = 16'h283;
#10;
address_ina = 252;
address_inb = 253;
data_ina = 16'h33e;
data_inb = 16'hfb68;
#10;
address_ina = 254;
address_inb = 255;
data_ina = 16'hfa10;
data_inb = 16'hffa2;
#10;
        wait(init_done);
        #30
        we = 0;
        // Start processing
         
		  #38000

        start = 0;



//        wait (wr_req);
//		  wait (!wr_req);
//		   rd_req = 1;
		  wait(done);
		  #20000
rd_req = 1;
        #70 
		  start = 1;
		 #80 
wait(rd_empty)
rd_req = 0;

$display("Finished the NTT test Number %d",test_num);
////Begin test number #33//////////////
rst = 1;

//#1000
start = 1;
mode = 1; //NTT 0 // INTT 1

// Reset for a few clock cycles

#1000

rst = 0;
test_num = test_num + 1;
#1000
we = 1;
address_ina = 0;
address_inb = 1;
data_ina = 16'h29f;
data_inb = 16'h1de;
#10;
address_ina = 2;
address_inb = 3;
data_ina = 16'h483;
data_inb = 16'hff55;
#10;
address_ina = 4;
address_inb = 5;
data_ina = 16'h311;
data_inb = 16'h317;
#10;
address_ina = 6;
address_inb = 7;
data_ina = 16'hfa0c;
data_inb = 16'hfc1d;
#10;
address_ina = 8;
address_inb = 9;
data_ina = 16'hfccf;
data_inb = 16'h208;
#10;
address_ina = 10;
address_inb = 11;
data_ina = 16'h1ea;
data_inb = 16'h605;
#10;
address_ina = 12;
address_inb = 13;
data_ina = 16'hfdea;
data_inb = 16'hfd99;
#10;
address_ina = 14;
address_inb = 15;
data_ina = 16'h17;
data_inb = 16'hfa79;
#10;
address_ina = 16;
address_inb = 17;
data_ina = 16'hfd32;
data_inb = 16'hfbc4;
#10;
address_ina = 18;
address_inb = 19;
data_ina = 16'hfd82;
data_inb = 16'hfabf;
#10;
address_ina = 20;
address_inb = 21;
data_ina = 16'h337;
data_inb = 16'hffac;
#10;
address_ina = 22;
address_inb = 23;
data_ina = 16'hfd8a;
data_inb = 16'ha3;
#10;
address_ina = 24;
address_inb = 25;
data_ina = 16'h537;
data_inb = 16'hffb7;
#10;
address_ina = 26;
address_inb = 27;
data_ina = 16'hfa5a;
data_inb = 16'h601;
#10;
address_ina = 28;
address_inb = 29;
data_ina = 16'h486;
data_inb = 16'hfa04;
#10;
address_ina = 30;
address_inb = 31;
data_ina = 16'hfa24;
data_inb = 16'h2cc;
#10;
address_ina = 32;
address_inb = 33;
data_ina = 16'h316;
data_inb = 16'hfa12;
#10;
address_ina = 34;
address_inb = 35;
data_ina = 16'hfb40;
data_inb = 16'h429;
#10;
address_ina = 36;
address_inb = 37;
data_ina = 16'h676;
data_inb = 16'hfc3f;
#10;
address_ina = 38;
address_inb = 39;
data_ina = 16'h501;
data_inb = 16'h647;
#10;
address_ina = 40;
address_inb = 41;
data_ina = 16'h506;
data_inb = 16'hfebe;
#10;
address_ina = 42;
address_inb = 43;
data_ina = 16'hfbdb;
data_inb = 16'h1c5;
#10;
address_ina = 44;
address_inb = 45;
data_ina = 16'hfb3d;
data_inb = 16'hfe85;
#10;
address_ina = 46;
address_inb = 47;
data_ina = 16'hff0e;
data_inb = 16'h2c9;
#10;
address_ina = 48;
address_inb = 49;
data_ina = 16'hfad8;
data_inb = 16'h54e;
#10;
address_ina = 50;
address_inb = 51;
data_ina = 16'h680;
data_inb = 16'h339;
#10;
address_ina = 52;
address_inb = 53;
data_ina = 16'h1cb;
data_inb = 16'hfdee;
#10;
address_ina = 54;
address_inb = 55;
data_ina = 16'h479;
data_inb = 16'hfec1;
#10;
address_ina = 56;
address_inb = 57;
data_ina = 16'hfe3a;
data_inb = 16'hfdd9;
#10;
address_ina = 58;
address_inb = 59;
data_ina = 16'hff0f;
data_inb = 16'h5fc;
#10;
address_ina = 60;
address_inb = 61;
data_ina = 16'hfa3b;
data_inb = 16'hfe71;
#10;
address_ina = 62;
address_inb = 63;
data_ina = 16'h2b0;
data_inb = 16'h9a;
#10;
address_ina = 64;
address_inb = 65;
data_ina = 16'hd6;
data_inb = 16'hfe9d;
#10;
address_ina = 66;
address_inb = 67;
data_ina = 16'h4e4;
data_inb = 16'h33a;
#10;
address_ina = 68;
address_inb = 69;
data_ina = 16'hfa28;
data_inb = 16'hfdd2;
#10;
address_ina = 70;
address_inb = 71;
data_ina = 16'hfe90;
data_inb = 16'h3a1;
#10;
address_ina = 72;
address_inb = 73;
data_ina = 16'hfdff;
data_inb = 16'h4ee;
#10;
address_ina = 74;
address_inb = 75;
data_ina = 16'hf9e0;
data_inb = 16'hf995;
#10;
address_ina = 76;
address_inb = 77;
data_ina = 16'hfa39;
data_inb = 16'h58c;
#10;
address_ina = 78;
address_inb = 79;
data_ina = 16'hfedb;
data_inb = 16'hf7;
#10;
address_ina = 80;
address_inb = 81;
data_ina = 16'hfc8f;
data_inb = 16'h64e;
#10;
address_ina = 82;
address_inb = 83;
data_ina = 16'h43c;
data_inb = 16'h432;
#10;
address_ina = 84;
address_inb = 85;
data_ina = 16'hfc89;
data_inb = 16'h18e;
#10;
address_ina = 86;
address_inb = 87;
data_ina = 16'h45f;
data_inb = 16'hfec9;
#10;
address_ina = 88;
address_inb = 89;
data_ina = 16'hffda;
data_inb = 16'hfe82;
#10;
address_ina = 90;
address_inb = 91;
data_ina = 16'hfb1d;
data_inb = 16'hfa2f;
#10;
address_ina = 92;
address_inb = 93;
data_ina = 16'h436;
data_inb = 16'h2da;
#10;
address_ina = 94;
address_inb = 95;
data_ina = 16'h4b1;
data_inb = 16'hfee5;
#10;
address_ina = 96;
address_inb = 97;
data_ina = 16'hfd91;
data_inb = 16'hfc53;
#10;
address_ina = 98;
address_inb = 99;
data_ina = 16'hfa75;
data_inb = 16'hfc7c;
#10;
address_ina = 100;
address_inb = 101;
data_ina = 16'hfe32;
data_inb = 16'h73;
#10;
address_ina = 102;
address_inb = 103;
data_ina = 16'h273;
data_inb = 16'h185;
#10;
address_ina = 104;
address_inb = 105;
data_ina = 16'h4c3;
data_inb = 16'h532;
#10;
address_ina = 106;
address_inb = 107;
data_ina = 16'h5ef;
data_inb = 16'h32a;
#10;
address_ina = 108;
address_inb = 109;
data_ina = 16'hfe25;
data_inb = 16'haf;
#10;
address_ina = 110;
address_inb = 111;
data_ina = 16'hfa97;
data_inb = 16'h199;
#10;
address_ina = 112;
address_inb = 113;
data_ina = 16'h66a;
data_inb = 16'hfd56;
#10;
address_ina = 114;
address_inb = 115;
data_ina = 16'h19;
data_inb = 16'h29e;
#10;
address_ina = 116;
address_inb = 117;
data_ina = 16'h187;
data_inb = 16'h52e;
#10;
address_ina = 118;
address_inb = 119;
data_ina = 16'h18c;
data_inb = 16'h440;
#10;
address_ina = 120;
address_inb = 121;
data_ina = 16'hfc29;
data_inb = 16'h56a;
#10;
address_ina = 122;
address_inb = 123;
data_ina = 16'hfd1c;
data_inb = 16'h183;
#10;
address_ina = 124;
address_inb = 125;
data_ina = 16'h413;
data_inb = 16'hfca8;
#10;
address_ina = 126;
address_inb = 127;
data_ina = 16'h39a;
data_inb = 16'hfac1;
#10;
address_ina = 128;
address_inb = 129;
data_ina = 16'h2a;
data_inb = 16'h5b1;
#10;
address_ina = 130;
address_inb = 131;
data_ina = 16'hfd63;
data_inb = 16'hfafc;
#10;
address_ina = 132;
address_inb = 133;
data_ina = 16'hfd5c;
data_inb = 16'h203;
#10;
address_ina = 134;
address_inb = 135;
data_ina = 16'hff77;
data_inb = 16'h390;
#10;
address_ina = 136;
address_inb = 137;
data_ina = 16'hfffb;
data_inb = 16'h63b;
#10;
address_ina = 138;
address_inb = 139;
data_ina = 16'h2ac;
data_inb = 16'h5f9;
#10;
address_ina = 140;
address_inb = 141;
data_ina = 16'hfd9a;
data_inb = 16'hfc20;
#10;
address_ina = 142;
address_inb = 143;
data_ina = 16'hfb29;
data_inb = 16'h2cc;
#10;
address_ina = 144;
address_inb = 145;
data_ina = 16'hfbc8;
data_inb = 16'hf9fd;
#10;
address_ina = 146;
address_inb = 147;
data_ina = 16'hffc0;
data_inb = 16'hfd96;
#10;
address_ina = 148;
address_inb = 149;
data_ina = 16'h298;
data_inb = 16'h31e;
#10;
address_ina = 150;
address_inb = 151;
data_ina = 16'hfc14;
data_inb = 16'h500;
#10;
address_ina = 152;
address_inb = 153;
data_ina = 16'hfc2f;
data_inb = 16'h2de;
#10;
address_ina = 154;
address_inb = 155;
data_ina = 16'h5c0;
data_inb = 16'h349;
#10;
address_ina = 156;
address_inb = 157;
data_ina = 16'h84;
data_inb = 16'hff80;
#10;
address_ina = 158;
address_inb = 159;
data_ina = 16'hfc22;
data_inb = 16'hfe18;
#10;
address_ina = 160;
address_inb = 161;
data_ina = 16'h51;
data_inb = 16'hbe;
#10;
address_ina = 162;
address_inb = 163;
data_ina = 16'hff04;
data_inb = 16'hfd2a;
#10;
address_ina = 164;
address_inb = 165;
data_ina = 16'hfb5d;
data_inb = 16'h51d;
#10;
address_ina = 166;
address_inb = 167;
data_ina = 16'hff4e;
data_inb = 16'hfc3a;
#10;
address_ina = 168;
address_inb = 169;
data_ina = 16'hac;
data_inb = 16'hfd45;
#10;
address_ina = 170;
address_inb = 171;
data_ina = 16'hfb84;
data_inb = 16'h39a;
#10;
address_ina = 172;
address_inb = 173;
data_ina = 16'hfa84;
data_inb = 16'hfc08;
#10;
address_ina = 174;
address_inb = 175;
data_ina = 16'h666;
data_inb = 16'h339;
#10;
address_ina = 176;
address_inb = 177;
data_ina = 16'hfd36;
data_inb = 16'hfc25;
#10;
address_ina = 178;
address_inb = 179;
data_ina = 16'h29a;
data_inb = 16'hff0c;
#10;
address_ina = 180;
address_inb = 181;
data_ina = 16'h42b;
data_inb = 16'hfe20;
#10;
address_ina = 182;
address_inb = 183;
data_ina = 16'h220;
data_inb = 16'hfa3d;
#10;
address_ina = 184;
address_inb = 185;
data_ina = 16'h56c;
data_inb = 16'h4df;
#10;
address_ina = 186;
address_inb = 187;
data_ina = 16'hfebf;
data_inb = 16'hca;
#10;
address_ina = 188;
address_inb = 189;
data_ina = 16'h298;
data_inb = 16'h5b7;
#10;
address_ina = 190;
address_inb = 191;
data_ina = 16'hfb66;
data_inb = 16'hfae2;
#10;
address_ina = 192;
address_inb = 193;
data_ina = 16'hff5b;
data_inb = 16'hfae7;
#10;
address_ina = 194;
address_inb = 195;
data_ina = 16'hfeda;
data_inb = 16'h1d4;
#10;
address_ina = 196;
address_inb = 197;
data_ina = 16'hfdda;
data_inb = 16'hfc0a;
#10;
address_ina = 198;
address_inb = 199;
data_ina = 16'h380;
data_inb = 16'hfa48;
#10;
address_ina = 200;
address_inb = 201;
data_ina = 16'hfdf1;
data_inb = 16'hfdfb;
#10;
address_ina = 202;
address_inb = 203;
data_ina = 16'hffca;
data_inb = 16'h445;
#10;
address_ina = 204;
address_inb = 205;
data_ina = 16'hfb53;
data_inb = 16'h54f;
#10;
address_ina = 206;
address_inb = 207;
data_ina = 16'hfa52;
data_inb = 16'hff5a;
#10;
address_ina = 208;
address_inb = 209;
data_ina = 16'hfdaf;
data_inb = 16'hfa4c;
#10;
address_ina = 210;
address_inb = 211;
data_ina = 16'hfa68;
data_inb = 16'hfe1a;
#10;
address_ina = 212;
address_inb = 213;
data_ina = 16'hfbdc;
data_inb = 16'hfc7d;
#10;
address_ina = 214;
address_inb = 215;
data_ina = 16'h5b1;
data_inb = 16'h3d3;
#10;
address_ina = 216;
address_inb = 217;
data_ina = 16'h282;
data_inb = 16'h5a3;
#10;
address_ina = 218;
address_inb = 219;
data_ina = 16'h230;
data_inb = 16'hfd43;
#10;
address_ina = 220;
address_inb = 221;
data_ina = 16'h4f4;
data_inb = 16'h35b;
#10;
address_ina = 222;
address_inb = 223;
data_ina = 16'h602;
data_inb = 16'h4aa;
#10;
address_ina = 224;
address_inb = 225;
data_ina = 16'h5ff;
data_inb = 16'h2de;
#10;
address_ina = 226;
address_inb = 227;
data_ina = 16'h370;
data_inb = 16'hfc92;
#10;
address_ina = 228;
address_inb = 229;
data_ina = 16'hfcc3;
data_inb = 16'h46d;
#10;
address_ina = 230;
address_inb = 231;
data_ina = 16'h106;
data_inb = 16'h2b6;
#10;
address_ina = 232;
address_inb = 233;
data_ina = 16'h152;
data_inb = 16'h2a9;
#10;
address_ina = 234;
address_inb = 235;
data_ina = 16'h3cf;
data_inb = 16'hfe12;
#10;
address_ina = 236;
address_inb = 237;
data_ina = 16'h380;
data_inb = 16'h520;
#10;
address_ina = 238;
address_inb = 239;
data_ina = 16'h558;
data_inb = 16'h72;
#10;
address_ina = 240;
address_inb = 241;
data_ina = 16'hf9db;
data_inb = 16'hfa36;
#10;
address_ina = 242;
address_inb = 243;
data_ina = 16'h9f;
data_inb = 16'h94;
#10;
address_ina = 244;
address_inb = 245;
data_ina = 16'hfa44;
data_inb = 16'h3d2;
#10;
address_ina = 246;
address_inb = 247;
data_ina = 16'h3fb;
data_inb = 16'hfa16;
#10;
address_ina = 248;
address_inb = 249;
data_ina = 16'hfce0;
data_inb = 16'hfc55;
#10;
address_ina = 250;
address_inb = 251;
data_ina = 16'hffbe;
data_inb = 16'h0;
#10;
address_ina = 252;
address_inb = 253;
data_ina = 16'hfe;
data_inb = 16'hface;
#10;
address_ina = 254;
address_inb = 255;
data_ina = 16'h674;
data_inb = 16'h2df;
#10;
        wait(init_done);
        #30
        we = 0;
        // Start processing
         
		  #38000

        start = 0;



//        wait (wr_req);
//		  wait (!wr_req);
//		   rd_req = 1;
		  wait(done);
		  #20000
rd_req = 1;
        #70 
		  start = 1;
		 #80 
wait(rd_empty)
rd_req = 0;

$display("Finished the NTT test Number %d",test_num);
////Begin test number #34//////////////
rst = 1;

//#1000
start = 1;
mode = 0; //NTT 0 // INTT 1

// Reset for a few clock cycles

#1000

rst = 0;
test_num = test_num + 1;
#1000
we = 1;
address_ina = 0;
address_inb = 1;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 2;
address_inb = 3;
data_ina = 16'h1;
data_inb = 16'h2;
#10;
address_ina = 4;
address_inb = 5;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 6;
address_inb = 7;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 8;
address_inb = 9;
data_ina = 16'hfffe;
data_inb = 16'h0;
#10;
address_ina = 10;
address_inb = 11;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 12;
address_inb = 13;
data_ina = 16'h1;
data_inb = 16'hfffe;
#10;
address_ina = 14;
address_inb = 15;
data_ina = 16'h2;
data_inb = 16'h2;
#10;
address_ina = 16;
address_inb = 17;
data_ina = 16'h2;
data_inb = 16'h2;
#10;
address_ina = 18;
address_inb = 19;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 20;
address_inb = 21;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 22;
address_inb = 23;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 24;
address_inb = 25;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 26;
address_inb = 27;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 28;
address_inb = 29;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 30;
address_inb = 31;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 32;
address_inb = 33;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 34;
address_inb = 35;
data_ina = 16'h1;
data_inb = 16'h2;
#10;
address_ina = 36;
address_inb = 37;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 38;
address_inb = 39;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 40;
address_inb = 41;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 42;
address_inb = 43;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 44;
address_inb = 45;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 46;
address_inb = 47;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 48;
address_inb = 49;
data_ina = 16'h0;
data_inb = 16'hfffe;
#10;
address_ina = 50;
address_inb = 51;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 52;
address_inb = 53;
data_ina = 16'hfffe;
data_inb = 16'h1;
#10;
address_ina = 54;
address_inb = 55;
data_ina = 16'h2;
data_inb = 16'h0;
#10;
address_ina = 56;
address_inb = 57;
data_ina = 16'h2;
data_inb = 16'hffff;
#10;
address_ina = 58;
address_inb = 59;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 60;
address_inb = 61;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 62;
address_inb = 63;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 64;
address_inb = 65;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 66;
address_inb = 67;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 68;
address_inb = 69;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 70;
address_inb = 71;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 72;
address_inb = 73;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 74;
address_inb = 75;
data_ina = 16'hffff;
data_inb = 16'h3;
#10;
address_ina = 76;
address_inb = 77;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 78;
address_inb = 79;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 80;
address_inb = 81;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 82;
address_inb = 83;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 84;
address_inb = 85;
data_ina = 16'h0;
data_inb = 16'h3;
#10;
address_ina = 86;
address_inb = 87;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 88;
address_inb = 89;
data_ina = 16'hffff;
data_inb = 16'h2;
#10;
address_ina = 90;
address_inb = 91;
data_ina = 16'hffff;
data_inb = 16'hfffe;
#10;
address_ina = 92;
address_inb = 93;
data_ina = 16'h2;
data_inb = 16'h2;
#10;
address_ina = 94;
address_inb = 95;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 96;
address_inb = 97;
data_ina = 16'h0;
data_inb = 16'h2;
#10;
address_ina = 98;
address_inb = 99;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 100;
address_inb = 101;
data_ina = 16'h2;
data_inb = 16'hffff;
#10;
address_ina = 102;
address_inb = 103;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 104;
address_inb = 105;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 106;
address_inb = 107;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 108;
address_inb = 109;
data_ina = 16'h1;
data_inb = 16'h2;
#10;
address_ina = 110;
address_inb = 111;
data_ina = 16'h0;
data_inb = 16'h2;
#10;
address_ina = 112;
address_inb = 113;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 114;
address_inb = 115;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 116;
address_inb = 117;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 118;
address_inb = 119;
data_ina = 16'hfffd;
data_inb = 16'hffff;
#10;
address_ina = 120;
address_inb = 121;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 122;
address_inb = 123;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 124;
address_inb = 125;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 126;
address_inb = 127;
data_ina = 16'h3;
data_inb = 16'h0;
#10;
address_ina = 128;
address_inb = 129;
data_ina = 16'h2;
data_inb = 16'h1;
#10;
address_ina = 130;
address_inb = 131;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 132;
address_inb = 133;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 134;
address_inb = 135;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 136;
address_inb = 137;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 138;
address_inb = 139;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 140;
address_inb = 141;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 142;
address_inb = 143;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 144;
address_inb = 145;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 146;
address_inb = 147;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 148;
address_inb = 149;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 150;
address_inb = 151;
data_ina = 16'h1;
data_inb = 16'hfffd;
#10;
address_ina = 152;
address_inb = 153;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 154;
address_inb = 155;
data_ina = 16'hfffe;
data_inb = 16'hfffe;
#10;
address_ina = 156;
address_inb = 157;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 158;
address_inb = 159;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 160;
address_inb = 161;
data_ina = 16'h0;
data_inb = 16'h2;
#10;
address_ina = 162;
address_inb = 163;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 164;
address_inb = 165;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 166;
address_inb = 167;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 168;
address_inb = 169;
data_ina = 16'h0;
data_inb = 16'hfffd;
#10;
address_ina = 170;
address_inb = 171;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 172;
address_inb = 173;
data_ina = 16'hfffe;
data_inb = 16'h1;
#10;
address_ina = 174;
address_inb = 175;
data_ina = 16'h0;
data_inb = 16'h2;
#10;
address_ina = 176;
address_inb = 177;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 178;
address_inb = 179;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 180;
address_inb = 181;
data_ina = 16'hfffe;
data_inb = 16'hfffe;
#10;
address_ina = 182;
address_inb = 183;
data_ina = 16'hffff;
data_inb = 16'hfffe;
#10;
address_ina = 184;
address_inb = 185;
data_ina = 16'h1;
data_inb = 16'hfffe;
#10;
address_ina = 186;
address_inb = 187;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 188;
address_inb = 189;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 190;
address_inb = 191;
data_ina = 16'h2;
data_inb = 16'h2;
#10;
address_ina = 192;
address_inb = 193;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 194;
address_inb = 195;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 196;
address_inb = 197;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 198;
address_inb = 199;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 200;
address_inb = 201;
data_ina = 16'h3;
data_inb = 16'h0;
#10;
address_ina = 202;
address_inb = 203;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 204;
address_inb = 205;
data_ina = 16'h2;
data_inb = 16'h0;
#10;
address_ina = 206;
address_inb = 207;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 208;
address_inb = 209;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 210;
address_inb = 211;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 212;
address_inb = 213;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 214;
address_inb = 215;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 216;
address_inb = 217;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 218;
address_inb = 219;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 220;
address_inb = 221;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 222;
address_inb = 223;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 224;
address_inb = 225;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 226;
address_inb = 227;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 228;
address_inb = 229;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 230;
address_inb = 231;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 232;
address_inb = 233;
data_ina = 16'hfffe;
data_inb = 16'h1;
#10;
address_ina = 234;
address_inb = 235;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 236;
address_inb = 237;
data_ina = 16'h0;
data_inb = 16'hfffe;
#10;
address_ina = 238;
address_inb = 239;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 240;
address_inb = 241;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 242;
address_inb = 243;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 244;
address_inb = 245;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 246;
address_inb = 247;
data_ina = 16'hfffd;
data_inb = 16'h1;
#10;
address_ina = 248;
address_inb = 249;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 250;
address_inb = 251;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 252;
address_inb = 253;
data_ina = 16'h2;
data_inb = 16'h0;
#10;
address_ina = 254;
address_inb = 255;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
        wait(init_done);
        #30
        we = 0;
        // Start processing
         
		  #38000

        start = 0;



//        wait (wr_req);
//		  wait (!wr_req);
//		   rd_req = 1;
		  wait(done);
		  #20000
rd_req = 1;
        #70 
		  start = 1;
		 #80 
wait(rd_empty)
rd_req = 0;

$display("Finished the NTT test Number %d",test_num);
////Begin test number #35//////////////
rst = 1;

//#1000
start = 1;
mode = 0; //NTT 0 // INTT 1

// Reset for a few clock cycles

#1000

rst = 0;
test_num = test_num + 1;
#1000
we = 1;
address_ina = 0;
address_inb = 1;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 2;
address_inb = 3;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 4;
address_inb = 5;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 6;
address_inb = 7;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 8;
address_inb = 9;
data_ina = 16'hffff;
data_inb = 16'h2;
#10;
address_ina = 10;
address_inb = 11;
data_ina = 16'h0;
data_inb = 16'h2;
#10;
address_ina = 12;
address_inb = 13;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 14;
address_inb = 15;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 16;
address_inb = 17;
data_ina = 16'h2;
data_inb = 16'hffff;
#10;
address_ina = 18;
address_inb = 19;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 20;
address_inb = 21;
data_ina = 16'h1;
data_inb = 16'hfffe;
#10;
address_ina = 22;
address_inb = 23;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 24;
address_inb = 25;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 26;
address_inb = 27;
data_ina = 16'h2;
data_inb = 16'h0;
#10;
address_ina = 28;
address_inb = 29;
data_ina = 16'hfffe;
data_inb = 16'hffff;
#10;
address_ina = 30;
address_inb = 31;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 32;
address_inb = 33;
data_ina = 16'h0;
data_inb = 16'h2;
#10;
address_ina = 34;
address_inb = 35;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 36;
address_inb = 37;
data_ina = 16'h0;
data_inb = 16'hfffe;
#10;
address_ina = 38;
address_inb = 39;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 40;
address_inb = 41;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 42;
address_inb = 43;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 44;
address_inb = 45;
data_ina = 16'h2;
data_inb = 16'hfffe;
#10;
address_ina = 46;
address_inb = 47;
data_ina = 16'h1;
data_inb = 16'h2;
#10;
address_ina = 48;
address_inb = 49;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 50;
address_inb = 51;
data_ina = 16'hfffe;
data_inb = 16'hffff;
#10;
address_ina = 52;
address_inb = 53;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 54;
address_inb = 55;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 56;
address_inb = 57;
data_ina = 16'h2;
data_inb = 16'h1;
#10;
address_ina = 58;
address_inb = 59;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 60;
address_inb = 61;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 62;
address_inb = 63;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 64;
address_inb = 65;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 66;
address_inb = 67;
data_ina = 16'h2;
data_inb = 16'hffff;
#10;
address_ina = 68;
address_inb = 69;
data_ina = 16'h0;
data_inb = 16'hfffe;
#10;
address_ina = 70;
address_inb = 71;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 72;
address_inb = 73;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 74;
address_inb = 75;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 76;
address_inb = 77;
data_ina = 16'hfffe;
data_inb = 16'h1;
#10;
address_ina = 78;
address_inb = 79;
data_ina = 16'h2;
data_inb = 16'h1;
#10;
address_ina = 80;
address_inb = 81;
data_ina = 16'h3;
data_inb = 16'hffff;
#10;
address_ina = 82;
address_inb = 83;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 84;
address_inb = 85;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 86;
address_inb = 87;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 88;
address_inb = 89;
data_ina = 16'hffff;
data_inb = 16'h2;
#10;
address_ina = 90;
address_inb = 91;
data_ina = 16'h2;
data_inb = 16'hffff;
#10;
address_ina = 92;
address_inb = 93;
data_ina = 16'h0;
data_inb = 16'h2;
#10;
address_ina = 94;
address_inb = 95;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 96;
address_inb = 97;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 98;
address_inb = 99;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 100;
address_inb = 101;
data_ina = 16'hffff;
data_inb = 16'h3;
#10;
address_ina = 102;
address_inb = 103;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 104;
address_inb = 105;
data_ina = 16'hffff;
data_inb = 16'h2;
#10;
address_ina = 106;
address_inb = 107;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 108;
address_inb = 109;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 110;
address_inb = 111;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 112;
address_inb = 113;
data_ina = 16'h1;
data_inb = 16'hfffe;
#10;
address_ina = 114;
address_inb = 115;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 116;
address_inb = 117;
data_ina = 16'h0;
data_inb = 16'h2;
#10;
address_ina = 118;
address_inb = 119;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 120;
address_inb = 121;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 122;
address_inb = 123;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 124;
address_inb = 125;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 126;
address_inb = 127;
data_ina = 16'h1;
data_inb = 16'h2;
#10;
address_ina = 128;
address_inb = 129;
data_ina = 16'h3;
data_inb = 16'h0;
#10;
address_ina = 130;
address_inb = 131;
data_ina = 16'h0;
data_inb = 16'hfffd;
#10;
address_ina = 132;
address_inb = 133;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 134;
address_inb = 135;
data_ina = 16'h0;
data_inb = 16'hfffe;
#10;
address_ina = 136;
address_inb = 137;
data_ina = 16'h0;
data_inb = 16'h2;
#10;
address_ina = 138;
address_inb = 139;
data_ina = 16'h0;
data_inb = 16'h2;
#10;
address_ina = 140;
address_inb = 141;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 142;
address_inb = 143;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 144;
address_inb = 145;
data_ina = 16'h2;
data_inb = 16'h1;
#10;
address_ina = 146;
address_inb = 147;
data_ina = 16'hfffe;
data_inb = 16'hffff;
#10;
address_ina = 148;
address_inb = 149;
data_ina = 16'h3;
data_inb = 16'h1;
#10;
address_ina = 150;
address_inb = 151;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 152;
address_inb = 153;
data_ina = 16'h0;
data_inb = 16'h2;
#10;
address_ina = 154;
address_inb = 155;
data_ina = 16'h1;
data_inb = 16'hfffe;
#10;
address_ina = 156;
address_inb = 157;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 158;
address_inb = 159;
data_ina = 16'hfffe;
data_inb = 16'h1;
#10;
address_ina = 160;
address_inb = 161;
data_ina = 16'h1;
data_inb = 16'h2;
#10;
address_ina = 162;
address_inb = 163;
data_ina = 16'h0;
data_inb = 16'h2;
#10;
address_ina = 164;
address_inb = 165;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 166;
address_inb = 167;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 168;
address_inb = 169;
data_ina = 16'hfffe;
data_inb = 16'h0;
#10;
address_ina = 170;
address_inb = 171;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 172;
address_inb = 173;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 174;
address_inb = 175;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 176;
address_inb = 177;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 178;
address_inb = 179;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 180;
address_inb = 181;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 182;
address_inb = 183;
data_ina = 16'h2;
data_inb = 16'h1;
#10;
address_ina = 184;
address_inb = 185;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 186;
address_inb = 187;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 188;
address_inb = 189;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 190;
address_inb = 191;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 192;
address_inb = 193;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 194;
address_inb = 195;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 196;
address_inb = 197;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 198;
address_inb = 199;
data_ina = 16'hffff;
data_inb = 16'hfffe;
#10;
address_ina = 200;
address_inb = 201;
data_ina = 16'hfffe;
data_inb = 16'hffff;
#10;
address_ina = 202;
address_inb = 203;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 204;
address_inb = 205;
data_ina = 16'h0;
data_inb = 16'h2;
#10;
address_ina = 206;
address_inb = 207;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 208;
address_inb = 209;
data_ina = 16'h0;
data_inb = 16'h2;
#10;
address_ina = 210;
address_inb = 211;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 212;
address_inb = 213;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 214;
address_inb = 215;
data_ina = 16'hffff;
data_inb = 16'hfffe;
#10;
address_ina = 216;
address_inb = 217;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 218;
address_inb = 219;
data_ina = 16'hfffe;
data_inb = 16'h1;
#10;
address_ina = 220;
address_inb = 221;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 222;
address_inb = 223;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 224;
address_inb = 225;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 226;
address_inb = 227;
data_ina = 16'h0;
data_inb = 16'hfffe;
#10;
address_ina = 228;
address_inb = 229;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 230;
address_inb = 231;
data_ina = 16'h3;
data_inb = 16'h1;
#10;
address_ina = 232;
address_inb = 233;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 234;
address_inb = 235;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 236;
address_inb = 237;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 238;
address_inb = 239;
data_ina = 16'hffff;
data_inb = 16'hfffe;
#10;
address_ina = 240;
address_inb = 241;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 242;
address_inb = 243;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 244;
address_inb = 245;
data_ina = 16'h2;
data_inb = 16'h0;
#10;
address_ina = 246;
address_inb = 247;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 248;
address_inb = 249;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 250;
address_inb = 251;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 252;
address_inb = 253;
data_ina = 16'hfffe;
data_inb = 16'h0;
#10;
address_ina = 254;
address_inb = 255;
data_ina = 16'h2;
data_inb = 16'h0;
#10;
        wait(init_done);
        #30
        we = 0;
        // Start processing
         
		  #38000

        start = 0;



//        wait (wr_req);
//		  wait (!wr_req);
//		   rd_req = 1;
		  wait(done);
		  #20000
rd_req = 1;
        #70 
		  start = 1;
		 #80 
wait(rd_empty)
rd_req = 0;

$display("Finished the NTT test Number %d",test_num);
////Begin test number #36//////////////
rst = 1;

//#1000
start = 1;
mode = 0; //NTT 0 // INTT 1

// Reset for a few clock cycles

#1000

rst = 0;
test_num = test_num + 1;
#1000
we = 1;
address_ina = 0;
address_inb = 1;
data_ina = 16'h2;
data_inb = 16'h0;
#10;
address_ina = 2;
address_inb = 3;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 4;
address_inb = 5;
data_ina = 16'h1;
data_inb = 16'hfffe;
#10;
address_ina = 6;
address_inb = 7;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 8;
address_inb = 9;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 10;
address_inb = 11;
data_ina = 16'h0;
data_inb = 16'h2;
#10;
address_ina = 12;
address_inb = 13;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 14;
address_inb = 15;
data_ina = 16'h1;
data_inb = 16'h3;
#10;
address_ina = 16;
address_inb = 17;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 18;
address_inb = 19;
data_ina = 16'hffff;
data_inb = 16'hfffe;
#10;
address_ina = 20;
address_inb = 21;
data_ina = 16'h2;
data_inb = 16'h0;
#10;
address_ina = 22;
address_inb = 23;
data_ina = 16'h2;
data_inb = 16'h1;
#10;
address_ina = 24;
address_inb = 25;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 26;
address_inb = 27;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 28;
address_inb = 29;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 30;
address_inb = 31;
data_ina = 16'h0;
data_inb = 16'hfffe;
#10;
address_ina = 32;
address_inb = 33;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 34;
address_inb = 35;
data_ina = 16'h2;
data_inb = 16'h1;
#10;
address_ina = 36;
address_inb = 37;
data_ina = 16'h2;
data_inb = 16'hffff;
#10;
address_ina = 38;
address_inb = 39;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 40;
address_inb = 41;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 42;
address_inb = 43;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 44;
address_inb = 45;
data_ina = 16'hfffe;
data_inb = 16'h1;
#10;
address_ina = 46;
address_inb = 47;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 48;
address_inb = 49;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 50;
address_inb = 51;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 52;
address_inb = 53;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 54;
address_inb = 55;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 56;
address_inb = 57;
data_ina = 16'h0;
data_inb = 16'hfffe;
#10;
address_ina = 58;
address_inb = 59;
data_ina = 16'h0;
data_inb = 16'h2;
#10;
address_ina = 60;
address_inb = 61;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 62;
address_inb = 63;
data_ina = 16'h0;
data_inb = 16'hfffe;
#10;
address_ina = 64;
address_inb = 65;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 66;
address_inb = 67;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 68;
address_inb = 69;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 70;
address_inb = 71;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 72;
address_inb = 73;
data_ina = 16'h2;
data_inb = 16'h1;
#10;
address_ina = 74;
address_inb = 75;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 76;
address_inb = 77;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 78;
address_inb = 79;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 80;
address_inb = 81;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 82;
address_inb = 83;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 84;
address_inb = 85;
data_ina = 16'h0;
data_inb = 16'h2;
#10;
address_ina = 86;
address_inb = 87;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 88;
address_inb = 89;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 90;
address_inb = 91;
data_ina = 16'h0;
data_inb = 16'hfffe;
#10;
address_ina = 92;
address_inb = 93;
data_ina = 16'h2;
data_inb = 16'h0;
#10;
address_ina = 94;
address_inb = 95;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 96;
address_inb = 97;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 98;
address_inb = 99;
data_ina = 16'h1;
data_inb = 16'h3;
#10;
address_ina = 100;
address_inb = 101;
data_ina = 16'h1;
data_inb = 16'hfffe;
#10;
address_ina = 102;
address_inb = 103;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 104;
address_inb = 105;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 106;
address_inb = 107;
data_ina = 16'hfffe;
data_inb = 16'h1;
#10;
address_ina = 108;
address_inb = 109;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 110;
address_inb = 111;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 112;
address_inb = 113;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 114;
address_inb = 115;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 116;
address_inb = 117;
data_ina = 16'h0;
data_inb = 16'h2;
#10;
address_ina = 118;
address_inb = 119;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 120;
address_inb = 121;
data_ina = 16'h0;
data_inb = 16'hfffe;
#10;
address_ina = 122;
address_inb = 123;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 124;
address_inb = 125;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 126;
address_inb = 127;
data_ina = 16'h2;
data_inb = 16'hffff;
#10;
address_ina = 128;
address_inb = 129;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 130;
address_inb = 131;
data_ina = 16'h0;
data_inb = 16'h2;
#10;
address_ina = 132;
address_inb = 133;
data_ina = 16'hfffe;
data_inb = 16'hfffd;
#10;
address_ina = 134;
address_inb = 135;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 136;
address_inb = 137;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 138;
address_inb = 139;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 140;
address_inb = 141;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 142;
address_inb = 143;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 144;
address_inb = 145;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 146;
address_inb = 147;
data_ina = 16'h2;
data_inb = 16'hffff;
#10;
address_ina = 148;
address_inb = 149;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 150;
address_inb = 151;
data_ina = 16'h0;
data_inb = 16'h2;
#10;
address_ina = 152;
address_inb = 153;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 154;
address_inb = 155;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 156;
address_inb = 157;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 158;
address_inb = 159;
data_ina = 16'h0;
data_inb = 16'h3;
#10;
address_ina = 160;
address_inb = 161;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 162;
address_inb = 163;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 164;
address_inb = 165;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 166;
address_inb = 167;
data_ina = 16'hfffe;
data_inb = 16'hffff;
#10;
address_ina = 168;
address_inb = 169;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 170;
address_inb = 171;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 172;
address_inb = 173;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 174;
address_inb = 175;
data_ina = 16'h2;
data_inb = 16'hfffe;
#10;
address_ina = 176;
address_inb = 177;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 178;
address_inb = 179;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 180;
address_inb = 181;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 182;
address_inb = 183;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 184;
address_inb = 185;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 186;
address_inb = 187;
data_ina = 16'hfffe;
data_inb = 16'h1;
#10;
address_ina = 188;
address_inb = 189;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 190;
address_inb = 191;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 192;
address_inb = 193;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 194;
address_inb = 195;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 196;
address_inb = 197;
data_ina = 16'h1;
data_inb = 16'hfffe;
#10;
address_ina = 198;
address_inb = 199;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 200;
address_inb = 201;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 202;
address_inb = 203;
data_ina = 16'h0;
data_inb = 16'hfffe;
#10;
address_ina = 204;
address_inb = 205;
data_ina = 16'hfffe;
data_inb = 16'hfffe;
#10;
address_ina = 206;
address_inb = 207;
data_ina = 16'hffff;
data_inb = 16'hfffe;
#10;
address_ina = 208;
address_inb = 209;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 210;
address_inb = 211;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 212;
address_inb = 213;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 214;
address_inb = 215;
data_ina = 16'hffff;
data_inb = 16'h3;
#10;
address_ina = 216;
address_inb = 217;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 218;
address_inb = 219;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 220;
address_inb = 221;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 222;
address_inb = 223;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 224;
address_inb = 225;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 226;
address_inb = 227;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 228;
address_inb = 229;
data_ina = 16'h2;
data_inb = 16'hffff;
#10;
address_ina = 230;
address_inb = 231;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 232;
address_inb = 233;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 234;
address_inb = 235;
data_ina = 16'h2;
data_inb = 16'hfffe;
#10;
address_ina = 236;
address_inb = 237;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 238;
address_inb = 239;
data_ina = 16'hfffe;
data_inb = 16'h1;
#10;
address_ina = 240;
address_inb = 241;
data_ina = 16'h2;
data_inb = 16'hffff;
#10;
address_ina = 242;
address_inb = 243;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 244;
address_inb = 245;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 246;
address_inb = 247;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 248;
address_inb = 249;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 250;
address_inb = 251;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 252;
address_inb = 253;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 254;
address_inb = 255;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
        wait(init_done);
        #30
        we = 0;
        // Start processing
         
		  #38000

        start = 0;



//        wait (wr_req);
//		  wait (!wr_req);
//		   rd_req = 1;
		  wait(done);
		  #20000
rd_req = 1;
        #70 
		  start = 1;
		 #80 
wait(rd_empty)
rd_req = 0;

$display("Finished the NTT test Number %d",test_num);
////Begin test number #37//////////////
rst = 1;

//#1000
start = 1;
mode = 0; //NTT 0 // INTT 1

// Reset for a few clock cycles

#1000

rst = 0;
test_num = test_num + 1;
#1000
we = 1;
address_ina = 0;
address_inb = 1;
data_ina = 16'hfffe;
data_inb = 16'h2;
#10;
address_ina = 2;
address_inb = 3;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 4;
address_inb = 5;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 6;
address_inb = 7;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 8;
address_inb = 9;
data_ina = 16'hfffd;
data_inb = 16'h1;
#10;
address_ina = 10;
address_inb = 11;
data_ina = 16'h1;
data_inb = 16'hfffe;
#10;
address_ina = 12;
address_inb = 13;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 14;
address_inb = 15;
data_ina = 16'hffff;
data_inb = 16'hfffe;
#10;
address_ina = 16;
address_inb = 17;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 18;
address_inb = 19;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 20;
address_inb = 21;
data_ina = 16'h0;
data_inb = 16'hfffd;
#10;
address_ina = 22;
address_inb = 23;
data_ina = 16'hfffe;
data_inb = 16'hffff;
#10;
address_ina = 24;
address_inb = 25;
data_ina = 16'h1;
data_inb = 16'hfffe;
#10;
address_ina = 26;
address_inb = 27;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 28;
address_inb = 29;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 30;
address_inb = 31;
data_ina = 16'hffff;
data_inb = 16'hfffe;
#10;
address_ina = 32;
address_inb = 33;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 34;
address_inb = 35;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 36;
address_inb = 37;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 38;
address_inb = 39;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 40;
address_inb = 41;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 42;
address_inb = 43;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 44;
address_inb = 45;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 46;
address_inb = 47;
data_ina = 16'h1;
data_inb = 16'hfffd;
#10;
address_ina = 48;
address_inb = 49;
data_ina = 16'h2;
data_inb = 16'h2;
#10;
address_ina = 50;
address_inb = 51;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 52;
address_inb = 53;
data_ina = 16'h0;
data_inb = 16'hfffe;
#10;
address_ina = 54;
address_inb = 55;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 56;
address_inb = 57;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 58;
address_inb = 59;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 60;
address_inb = 61;
data_ina = 16'h1;
data_inb = 16'hfffe;
#10;
address_ina = 62;
address_inb = 63;
data_ina = 16'h1;
data_inb = 16'hfffd;
#10;
address_ina = 64;
address_inb = 65;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 66;
address_inb = 67;
data_ina = 16'h2;
data_inb = 16'hfffe;
#10;
address_ina = 68;
address_inb = 69;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 70;
address_inb = 71;
data_ina = 16'hfffe;
data_inb = 16'hffff;
#10;
address_ina = 72;
address_inb = 73;
data_ina = 16'h0;
data_inb = 16'hfffe;
#10;
address_ina = 74;
address_inb = 75;
data_ina = 16'hfffe;
data_inb = 16'h2;
#10;
address_ina = 76;
address_inb = 77;
data_ina = 16'h2;
data_inb = 16'hffff;
#10;
address_ina = 78;
address_inb = 79;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 80;
address_inb = 81;
data_ina = 16'hffff;
data_inb = 16'h2;
#10;
address_ina = 82;
address_inb = 83;
data_ina = 16'h0;
data_inb = 16'hfffe;
#10;
address_ina = 84;
address_inb = 85;
data_ina = 16'h2;
data_inb = 16'h1;
#10;
address_ina = 86;
address_inb = 87;
data_ina = 16'hffff;
data_inb = 16'h2;
#10;
address_ina = 88;
address_inb = 89;
data_ina = 16'hfffe;
data_inb = 16'h1;
#10;
address_ina = 90;
address_inb = 91;
data_ina = 16'h2;
data_inb = 16'hfffe;
#10;
address_ina = 92;
address_inb = 93;
data_ina = 16'hfffe;
data_inb = 16'h2;
#10;
address_ina = 94;
address_inb = 95;
data_ina = 16'h0;
data_inb = 16'hfffe;
#10;
address_ina = 96;
address_inb = 97;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 98;
address_inb = 99;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 100;
address_inb = 101;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 102;
address_inb = 103;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 104;
address_inb = 105;
data_ina = 16'h0;
data_inb = 16'hfffe;
#10;
address_ina = 106;
address_inb = 107;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 108;
address_inb = 109;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 110;
address_inb = 111;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 112;
address_inb = 113;
data_ina = 16'h0;
data_inb = 16'hfffe;
#10;
address_ina = 114;
address_inb = 115;
data_ina = 16'hfffe;
data_inb = 16'h2;
#10;
address_ina = 116;
address_inb = 117;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 118;
address_inb = 119;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 120;
address_inb = 121;
data_ina = 16'h3;
data_inb = 16'h0;
#10;
address_ina = 122;
address_inb = 123;
data_ina = 16'hfffd;
data_inb = 16'h0;
#10;
address_ina = 124;
address_inb = 125;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 126;
address_inb = 127;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 128;
address_inb = 129;
data_ina = 16'hfffe;
data_inb = 16'h0;
#10;
address_ina = 130;
address_inb = 131;
data_ina = 16'h2;
data_inb = 16'h0;
#10;
address_ina = 132;
address_inb = 133;
data_ina = 16'hffff;
data_inb = 16'hfffe;
#10;
address_ina = 134;
address_inb = 135;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 136;
address_inb = 137;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 138;
address_inb = 139;
data_ina = 16'h2;
data_inb = 16'h0;
#10;
address_ina = 140;
address_inb = 141;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 142;
address_inb = 143;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 144;
address_inb = 145;
data_ina = 16'h1;
data_inb = 16'h2;
#10;
address_ina = 146;
address_inb = 147;
data_ina = 16'hfffe;
data_inb = 16'h2;
#10;
address_ina = 148;
address_inb = 149;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 150;
address_inb = 151;
data_ina = 16'hfffe;
data_inb = 16'h2;
#10;
address_ina = 152;
address_inb = 153;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 154;
address_inb = 155;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 156;
address_inb = 157;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 158;
address_inb = 159;
data_ina = 16'h3;
data_inb = 16'hffff;
#10;
address_ina = 160;
address_inb = 161;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 162;
address_inb = 163;
data_ina = 16'h2;
data_inb = 16'h2;
#10;
address_ina = 164;
address_inb = 165;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 166;
address_inb = 167;
data_ina = 16'h0;
data_inb = 16'h2;
#10;
address_ina = 168;
address_inb = 169;
data_ina = 16'hfffe;
data_inb = 16'h0;
#10;
address_ina = 170;
address_inb = 171;
data_ina = 16'h2;
data_inb = 16'hffff;
#10;
address_ina = 172;
address_inb = 173;
data_ina = 16'h2;
data_inb = 16'h0;
#10;
address_ina = 174;
address_inb = 175;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 176;
address_inb = 177;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 178;
address_inb = 179;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 180;
address_inb = 181;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 182;
address_inb = 183;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 184;
address_inb = 185;
data_ina = 16'h1;
data_inb = 16'h2;
#10;
address_ina = 186;
address_inb = 187;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 188;
address_inb = 189;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 190;
address_inb = 191;
data_ina = 16'hffff;
data_inb = 16'h3;
#10;
address_ina = 192;
address_inb = 193;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 194;
address_inb = 195;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 196;
address_inb = 197;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 198;
address_inb = 199;
data_ina = 16'h2;
data_inb = 16'h0;
#10;
address_ina = 200;
address_inb = 201;
data_ina = 16'h1;
data_inb = 16'h3;
#10;
address_ina = 202;
address_inb = 203;
data_ina = 16'h0;
data_inb = 16'hfffd;
#10;
address_ina = 204;
address_inb = 205;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 206;
address_inb = 207;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 208;
address_inb = 209;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 210;
address_inb = 211;
data_ina = 16'h0;
data_inb = 16'hfffe;
#10;
address_ina = 212;
address_inb = 213;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 214;
address_inb = 215;
data_ina = 16'hfffe;
data_inb = 16'h1;
#10;
address_ina = 216;
address_inb = 217;
data_ina = 16'h3;
data_inb = 16'h1;
#10;
address_ina = 218;
address_inb = 219;
data_ina = 16'hfffe;
data_inb = 16'hffff;
#10;
address_ina = 220;
address_inb = 221;
data_ina = 16'hffff;
data_inb = 16'hfffe;
#10;
address_ina = 222;
address_inb = 223;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 224;
address_inb = 225;
data_ina = 16'h2;
data_inb = 16'h0;
#10;
address_ina = 226;
address_inb = 227;
data_ina = 16'hfffe;
data_inb = 16'h0;
#10;
address_ina = 228;
address_inb = 229;
data_ina = 16'hfffe;
data_inb = 16'h2;
#10;
address_ina = 230;
address_inb = 231;
data_ina = 16'h2;
data_inb = 16'hffff;
#10;
address_ina = 232;
address_inb = 233;
data_ina = 16'h2;
data_inb = 16'h1;
#10;
address_ina = 234;
address_inb = 235;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 236;
address_inb = 237;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 238;
address_inb = 239;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 240;
address_inb = 241;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 242;
address_inb = 243;
data_ina = 16'h2;
data_inb = 16'h1;
#10;
address_ina = 244;
address_inb = 245;
data_ina = 16'h1;
data_inb = 16'hfffd;
#10;
address_ina = 246;
address_inb = 247;
data_ina = 16'hfffe;
data_inb = 16'h1;
#10;
address_ina = 248;
address_inb = 249;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 250;
address_inb = 251;
data_ina = 16'hffff;
data_inb = 16'hfffe;
#10;
address_ina = 252;
address_inb = 253;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 254;
address_inb = 255;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
        wait(init_done);
        #30
        we = 0;
        // Start processing
         
		  #38000

        start = 0;



//        wait (wr_req);
//		  wait (!wr_req);
//		   rd_req = 1;
		  wait(done);
		  #20000
rd_req = 1;
        #70 
		  start = 1;
		 #80 
wait(rd_empty)
rd_req = 0;

$display("Finished the NTT test Number %d",test_num);
////Begin test number #38//////////////
rst = 1;

//#1000
start = 1;
mode = 0; //NTT 0 // INTT 1

// Reset for a few clock cycles

#1000

rst = 0;
test_num = test_num + 1;
#1000
we = 1;
address_ina = 0;
address_inb = 1;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 2;
address_inb = 3;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 4;
address_inb = 5;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 6;
address_inb = 7;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 8;
address_inb = 9;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 10;
address_inb = 11;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 12;
address_inb = 13;
data_ina = 16'h0;
data_inb = 16'h2;
#10;
address_ina = 14;
address_inb = 15;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 16;
address_inb = 17;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 18;
address_inb = 19;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 20;
address_inb = 21;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 22;
address_inb = 23;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 24;
address_inb = 25;
data_ina = 16'hfffe;
data_inb = 16'hfffe;
#10;
address_ina = 26;
address_inb = 27;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 28;
address_inb = 29;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 30;
address_inb = 31;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 32;
address_inb = 33;
data_ina = 16'h0;
data_inb = 16'h2;
#10;
address_ina = 34;
address_inb = 35;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 36;
address_inb = 37;
data_ina = 16'h1;
data_inb = 16'hfffe;
#10;
address_ina = 38;
address_inb = 39;
data_ina = 16'h2;
data_inb = 16'hfffe;
#10;
address_ina = 40;
address_inb = 41;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 42;
address_inb = 43;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 44;
address_inb = 45;
data_ina = 16'h0;
data_inb = 16'h2;
#10;
address_ina = 46;
address_inb = 47;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 48;
address_inb = 49;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 50;
address_inb = 51;
data_ina = 16'hfffe;
data_inb = 16'h0;
#10;
address_ina = 52;
address_inb = 53;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 54;
address_inb = 55;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 56;
address_inb = 57;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 58;
address_inb = 59;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 60;
address_inb = 61;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 62;
address_inb = 63;
data_ina = 16'h2;
data_inb = 16'hffff;
#10;
address_ina = 64;
address_inb = 65;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 66;
address_inb = 67;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 68;
address_inb = 69;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 70;
address_inb = 71;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 72;
address_inb = 73;
data_ina = 16'hffff;
data_inb = 16'hfffe;
#10;
address_ina = 74;
address_inb = 75;
data_ina = 16'h2;
data_inb = 16'h0;
#10;
address_ina = 76;
address_inb = 77;
data_ina = 16'hffff;
data_inb = 16'h2;
#10;
address_ina = 78;
address_inb = 79;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 80;
address_inb = 81;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 82;
address_inb = 83;
data_ina = 16'h2;
data_inb = 16'h0;
#10;
address_ina = 84;
address_inb = 85;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 86;
address_inb = 87;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 88;
address_inb = 89;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 90;
address_inb = 91;
data_ina = 16'hffff;
data_inb = 16'hfffe;
#10;
address_ina = 92;
address_inb = 93;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 94;
address_inb = 95;
data_ina = 16'h2;
data_inb = 16'h1;
#10;
address_ina = 96;
address_inb = 97;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 98;
address_inb = 99;
data_ina = 16'h0;
data_inb = 16'h2;
#10;
address_ina = 100;
address_inb = 101;
data_ina = 16'h0;
data_inb = 16'hfffe;
#10;
address_ina = 102;
address_inb = 103;
data_ina = 16'h2;
data_inb = 16'h0;
#10;
address_ina = 104;
address_inb = 105;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 106;
address_inb = 107;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 108;
address_inb = 109;
data_ina = 16'hfffe;
data_inb = 16'hffff;
#10;
address_ina = 110;
address_inb = 111;
data_ina = 16'hfffd;
data_inb = 16'h1;
#10;
address_ina = 112;
address_inb = 113;
data_ina = 16'h0;
data_inb = 16'hfffe;
#10;
address_ina = 114;
address_inb = 115;
data_ina = 16'hfffe;
data_inb = 16'hfffe;
#10;
address_ina = 116;
address_inb = 117;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 118;
address_inb = 119;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 120;
address_inb = 121;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 122;
address_inb = 123;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 124;
address_inb = 125;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 126;
address_inb = 127;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 128;
address_inb = 129;
data_ina = 16'h2;
data_inb = 16'hfffd;
#10;
address_ina = 130;
address_inb = 131;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 132;
address_inb = 133;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 134;
address_inb = 135;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 136;
address_inb = 137;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 138;
address_inb = 139;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 140;
address_inb = 141;
data_ina = 16'h0;
data_inb = 16'h2;
#10;
address_ina = 142;
address_inb = 143;
data_ina = 16'hfffd;
data_inb = 16'h0;
#10;
address_ina = 144;
address_inb = 145;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 146;
address_inb = 147;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 148;
address_inb = 149;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 150;
address_inb = 151;
data_ina = 16'h2;
data_inb = 16'h0;
#10;
address_ina = 152;
address_inb = 153;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 154;
address_inb = 155;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 156;
address_inb = 157;
data_ina = 16'h0;
data_inb = 16'hfffe;
#10;
address_ina = 158;
address_inb = 159;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 160;
address_inb = 161;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 162;
address_inb = 163;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 164;
address_inb = 165;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 166;
address_inb = 167;
data_ina = 16'h2;
data_inb = 16'h0;
#10;
address_ina = 168;
address_inb = 169;
data_ina = 16'hffff;
data_inb = 16'h2;
#10;
address_ina = 170;
address_inb = 171;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 172;
address_inb = 173;
data_ina = 16'hffff;
data_inb = 16'hfffe;
#10;
address_ina = 174;
address_inb = 175;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 176;
address_inb = 177;
data_ina = 16'h2;
data_inb = 16'h2;
#10;
address_ina = 178;
address_inb = 179;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 180;
address_inb = 181;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 182;
address_inb = 183;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 184;
address_inb = 185;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 186;
address_inb = 187;
data_ina = 16'h3;
data_inb = 16'h0;
#10;
address_ina = 188;
address_inb = 189;
data_ina = 16'hfffe;
data_inb = 16'h3;
#10;
address_ina = 190;
address_inb = 191;
data_ina = 16'h0;
data_inb = 16'h2;
#10;
address_ina = 192;
address_inb = 193;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 194;
address_inb = 195;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 196;
address_inb = 197;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 198;
address_inb = 199;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 200;
address_inb = 201;
data_ina = 16'hfffe;
data_inb = 16'h1;
#10;
address_ina = 202;
address_inb = 203;
data_ina = 16'h0;
data_inb = 16'h2;
#10;
address_ina = 204;
address_inb = 205;
data_ina = 16'h0;
data_inb = 16'hfffe;
#10;
address_ina = 206;
address_inb = 207;
data_ina = 16'h2;
data_inb = 16'h0;
#10;
address_ina = 208;
address_inb = 209;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 210;
address_inb = 211;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 212;
address_inb = 213;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 214;
address_inb = 215;
data_ina = 16'hfffd;
data_inb = 16'hffff;
#10;
address_ina = 216;
address_inb = 217;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 218;
address_inb = 219;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 220;
address_inb = 221;
data_ina = 16'hfffe;
data_inb = 16'h0;
#10;
address_ina = 222;
address_inb = 223;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 224;
address_inb = 225;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 226;
address_inb = 227;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 228;
address_inb = 229;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 230;
address_inb = 231;
data_ina = 16'h2;
data_inb = 16'h1;
#10;
address_ina = 232;
address_inb = 233;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 234;
address_inb = 235;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 236;
address_inb = 237;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 238;
address_inb = 239;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 240;
address_inb = 241;
data_ina = 16'h0;
data_inb = 16'hfffe;
#10;
address_ina = 242;
address_inb = 243;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 244;
address_inb = 245;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 246;
address_inb = 247;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 248;
address_inb = 249;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 250;
address_inb = 251;
data_ina = 16'h2;
data_inb = 16'h3;
#10;
address_ina = 252;
address_inb = 253;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 254;
address_inb = 255;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
        wait(init_done);
        #30
        we = 0;
        // Start processing
         
		  #38000

        start = 0;



//        wait (wr_req);
//		  wait (!wr_req);
//		   rd_req = 1;
		  wait(done);
		  #20000
rd_req = 1;
        #70 
		  start = 1;
		 #80 
wait(rd_empty)
rd_req = 0;

$display("Finished the NTT test Number %d",test_num);
////Begin test number #39//////////////
rst = 1;

//#1000
start = 1;
mode = 0; //NTT 0 // INTT 1

// Reset for a few clock cycles

#1000

rst = 0;
test_num = test_num + 1;
#1000
we = 1;
address_ina = 0;
address_inb = 1;
data_ina = 16'h1;
data_inb = 16'hfffe;
#10;
address_ina = 2;
address_inb = 3;
data_ina = 16'h2;
data_inb = 16'hffff;
#10;
address_ina = 4;
address_inb = 5;
data_ina = 16'hfffe;
data_inb = 16'hffff;
#10;
address_ina = 6;
address_inb = 7;
data_ina = 16'h2;
data_inb = 16'h0;
#10;
address_ina = 8;
address_inb = 9;
data_ina = 16'hfffe;
data_inb = 16'h0;
#10;
address_ina = 10;
address_inb = 11;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 12;
address_inb = 13;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 14;
address_inb = 15;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 16;
address_inb = 17;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 18;
address_inb = 19;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 20;
address_inb = 21;
data_ina = 16'hfffe;
data_inb = 16'h1;
#10;
address_ina = 22;
address_inb = 23;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 24;
address_inb = 25;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 26;
address_inb = 27;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 28;
address_inb = 29;
data_ina = 16'hffff;
data_inb = 16'hfffe;
#10;
address_ina = 30;
address_inb = 31;
data_ina = 16'h2;
data_inb = 16'hfffe;
#10;
address_ina = 32;
address_inb = 33;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 34;
address_inb = 35;
data_ina = 16'h2;
data_inb = 16'h0;
#10;
address_ina = 36;
address_inb = 37;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 38;
address_inb = 39;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 40;
address_inb = 41;
data_ina = 16'h2;
data_inb = 16'h3;
#10;
address_ina = 42;
address_inb = 43;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 44;
address_inb = 45;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 46;
address_inb = 47;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 48;
address_inb = 49;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 50;
address_inb = 51;
data_ina = 16'h1;
data_inb = 16'hfffe;
#10;
address_ina = 52;
address_inb = 53;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 54;
address_inb = 55;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 56;
address_inb = 57;
data_ina = 16'hfffe;
data_inb = 16'hffff;
#10;
address_ina = 58;
address_inb = 59;
data_ina = 16'hffff;
data_inb = 16'h2;
#10;
address_ina = 60;
address_inb = 61;
data_ina = 16'hfffe;
data_inb = 16'h0;
#10;
address_ina = 62;
address_inb = 63;
data_ina = 16'hffff;
data_inb = 16'h2;
#10;
address_ina = 64;
address_inb = 65;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 66;
address_inb = 67;
data_ina = 16'h2;
data_inb = 16'h0;
#10;
address_ina = 68;
address_inb = 69;
data_ina = 16'h0;
data_inb = 16'hfffe;
#10;
address_ina = 70;
address_inb = 71;
data_ina = 16'h1;
data_inb = 16'h2;
#10;
address_ina = 72;
address_inb = 73;
data_ina = 16'hfffd;
data_inb = 16'h0;
#10;
address_ina = 74;
address_inb = 75;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 76;
address_inb = 77;
data_ina = 16'hfffe;
data_inb = 16'h0;
#10;
address_ina = 78;
address_inb = 79;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 80;
address_inb = 81;
data_ina = 16'hfffe;
data_inb = 16'hffff;
#10;
address_ina = 82;
address_inb = 83;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 84;
address_inb = 85;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 86;
address_inb = 87;
data_ina = 16'hfffe;
data_inb = 16'h2;
#10;
address_ina = 88;
address_inb = 89;
data_ina = 16'hfffd;
data_inb = 16'h1;
#10;
address_ina = 90;
address_inb = 91;
data_ina = 16'h0;
data_inb = 16'hfffe;
#10;
address_ina = 92;
address_inb = 93;
data_ina = 16'h0;
data_inb = 16'h3;
#10;
address_ina = 94;
address_inb = 95;
data_ina = 16'hfffe;
data_inb = 16'h2;
#10;
address_ina = 96;
address_inb = 97;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 98;
address_inb = 99;
data_ina = 16'hfffe;
data_inb = 16'hfffe;
#10;
address_ina = 100;
address_inb = 101;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 102;
address_inb = 103;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 104;
address_inb = 105;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 106;
address_inb = 107;
data_ina = 16'h0;
data_inb = 16'h3;
#10;
address_ina = 108;
address_inb = 109;
data_ina = 16'h0;
data_inb = 16'hfffe;
#10;
address_ina = 110;
address_inb = 111;
data_ina = 16'h1;
data_inb = 16'hfffe;
#10;
address_ina = 112;
address_inb = 113;
data_ina = 16'h2;
data_inb = 16'h0;
#10;
address_ina = 114;
address_inb = 115;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 116;
address_inb = 117;
data_ina = 16'h0;
data_inb = 16'h3;
#10;
address_ina = 118;
address_inb = 119;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 120;
address_inb = 121;
data_ina = 16'hffff;
data_inb = 16'hfffe;
#10;
address_ina = 122;
address_inb = 123;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 124;
address_inb = 125;
data_ina = 16'hfffe;
data_inb = 16'hffff;
#10;
address_ina = 126;
address_inb = 127;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 128;
address_inb = 129;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 130;
address_inb = 131;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 132;
address_inb = 133;
data_ina = 16'h1;
data_inb = 16'hfffe;
#10;
address_ina = 134;
address_inb = 135;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 136;
address_inb = 137;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 138;
address_inb = 139;
data_ina = 16'hfffe;
data_inb = 16'h0;
#10;
address_ina = 140;
address_inb = 141;
data_ina = 16'h1;
data_inb = 16'hfffe;
#10;
address_ina = 142;
address_inb = 143;
data_ina = 16'hffff;
data_inb = 16'h2;
#10;
address_ina = 144;
address_inb = 145;
data_ina = 16'h2;
data_inb = 16'h0;
#10;
address_ina = 146;
address_inb = 147;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 148;
address_inb = 149;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 150;
address_inb = 151;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 152;
address_inb = 153;
data_ina = 16'hffff;
data_inb = 16'h2;
#10;
address_ina = 154;
address_inb = 155;
data_ina = 16'h0;
data_inb = 16'h2;
#10;
address_ina = 156;
address_inb = 157;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 158;
address_inb = 159;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 160;
address_inb = 161;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 162;
address_inb = 163;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 164;
address_inb = 165;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 166;
address_inb = 167;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 168;
address_inb = 169;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 170;
address_inb = 171;
data_ina = 16'h2;
data_inb = 16'h0;
#10;
address_ina = 172;
address_inb = 173;
data_ina = 16'hffff;
data_inb = 16'hfffe;
#10;
address_ina = 174;
address_inb = 175;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 176;
address_inb = 177;
data_ina = 16'h2;
data_inb = 16'h0;
#10;
address_ina = 178;
address_inb = 179;
data_ina = 16'h2;
data_inb = 16'h1;
#10;
address_ina = 180;
address_inb = 181;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 182;
address_inb = 183;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 184;
address_inb = 185;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 186;
address_inb = 187;
data_ina = 16'hffff;
data_inb = 16'h2;
#10;
address_ina = 188;
address_inb = 189;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 190;
address_inb = 191;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 192;
address_inb = 193;
data_ina = 16'h0;
data_inb = 16'hfffe;
#10;
address_ina = 194;
address_inb = 195;
data_ina = 16'h1;
data_inb = 16'h2;
#10;
address_ina = 196;
address_inb = 197;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 198;
address_inb = 199;
data_ina = 16'hffff;
data_inb = 16'hfffe;
#10;
address_ina = 200;
address_inb = 201;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 202;
address_inb = 203;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 204;
address_inb = 205;
data_ina = 16'h0;
data_inb = 16'h3;
#10;
address_ina = 206;
address_inb = 207;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 208;
address_inb = 209;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 210;
address_inb = 211;
data_ina = 16'h2;
data_inb = 16'h2;
#10;
address_ina = 212;
address_inb = 213;
data_ina = 16'h2;
data_inb = 16'h1;
#10;
address_ina = 214;
address_inb = 215;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 216;
address_inb = 217;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 218;
address_inb = 219;
data_ina = 16'hfffe;
data_inb = 16'h0;
#10;
address_ina = 220;
address_inb = 221;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 222;
address_inb = 223;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 224;
address_inb = 225;
data_ina = 16'h2;
data_inb = 16'h0;
#10;
address_ina = 226;
address_inb = 227;
data_ina = 16'h3;
data_inb = 16'h0;
#10;
address_ina = 228;
address_inb = 229;
data_ina = 16'hfffe;
data_inb = 16'h1;
#10;
address_ina = 230;
address_inb = 231;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 232;
address_inb = 233;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 234;
address_inb = 235;
data_ina = 16'hffff;
data_inb = 16'hfffe;
#10;
address_ina = 236;
address_inb = 237;
data_ina = 16'hffff;
data_inb = 16'hfffe;
#10;
address_ina = 238;
address_inb = 239;
data_ina = 16'hffff;
data_inb = 16'hfffe;
#10;
address_ina = 240;
address_inb = 241;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 242;
address_inb = 243;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 244;
address_inb = 245;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 246;
address_inb = 247;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 248;
address_inb = 249;
data_ina = 16'hfffe;
data_inb = 16'h2;
#10;
address_ina = 250;
address_inb = 251;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 252;
address_inb = 253;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 254;
address_inb = 255;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
        wait(init_done);
        #30
        we = 0;
        // Start processing
         
		  #38000

        start = 0;



//        wait (wr_req);
//		  wait (!wr_req);
//		   rd_req = 1;
		  wait(done);
		  #20000
rd_req = 1;
        #70 
		  start = 1;
		 #80 
wait(rd_empty)
rd_req = 0;

$display("Finished the NTT test Number %d",test_num);
////Begin test number #40//////////////
rst = 1;

//#1000
start = 1;
mode = 1; //NTT 0 // INTT 1

// Reset for a few clock cycles

#1000

rst = 0;
test_num = test_num + 1;
#1000
we = 1;
address_ina = 0;
address_inb = 1;
data_ina = 16'hf9e0;
data_inb = 16'hfa0e;
#10;
address_ina = 2;
address_inb = 3;
data_ina = 16'h43;
data_inb = 16'hfb61;
#10;
address_ina = 4;
address_inb = 5;
data_ina = 16'h2f7;
data_inb = 16'hff7d;
#10;
address_ina = 6;
address_inb = 7;
data_ina = 16'h5c6;
data_inb = 16'h29d;
#10;
address_ina = 8;
address_inb = 9;
data_ina = 16'hfc52;
data_inb = 16'hff76;
#10;
address_ina = 10;
address_inb = 11;
data_ina = 16'h4fa;
data_inb = 16'h2ef;
#10;
address_ina = 12;
address_inb = 13;
data_ina = 16'h555;
data_inb = 16'h4fd;
#10;
address_ina = 14;
address_inb = 15;
data_ina = 16'hfdc3;
data_inb = 16'hfec1;
#10;
address_ina = 16;
address_inb = 17;
data_ina = 16'h54d;
data_inb = 16'h5d0;
#10;
address_ina = 18;
address_inb = 19;
data_ina = 16'h454;
data_inb = 16'hff6d;
#10;
address_ina = 20;
address_inb = 21;
data_ina = 16'hfb53;
data_inb = 16'hffd9;
#10;
address_ina = 22;
address_inb = 23;
data_ina = 16'he9;
data_inb = 16'hfce4;
#10;
address_ina = 24;
address_inb = 25;
data_ina = 16'hfb46;
data_inb = 16'h65d;
#10;
address_ina = 26;
address_inb = 27;
data_ina = 16'hffcf;
data_inb = 16'hfe85;
#10;
address_ina = 28;
address_inb = 29;
data_ina = 16'h174;
data_inb = 16'h15a;
#10;
address_ina = 30;
address_inb = 31;
data_ina = 16'h129;
data_inb = 16'hfaa8;
#10;
address_ina = 32;
address_inb = 33;
data_ina = 16'hfe3e;
data_inb = 16'h72;
#10;
address_ina = 34;
address_inb = 35;
data_ina = 16'hfb02;
data_inb = 16'h3e3;
#10;
address_ina = 36;
address_inb = 37;
data_ina = 16'h30e;
data_inb = 16'h10a;
#10;
address_ina = 38;
address_inb = 39;
data_ina = 16'hfbcc;
data_inb = 16'hfdc1;
#10;
address_ina = 40;
address_inb = 41;
data_ina = 16'hff11;
data_inb = 16'h5ad;
#10;
address_ina = 42;
address_inb = 43;
data_ina = 16'h676;
data_inb = 16'hfb16;
#10;
address_ina = 44;
address_inb = 45;
data_ina = 16'haa;
data_inb = 16'hfed1;
#10;
address_ina = 46;
address_inb = 47;
data_ina = 16'hfcdc;
data_inb = 16'hfbc6;
#10;
address_ina = 48;
address_inb = 49;
data_ina = 16'h43f;
data_inb = 16'hfb1f;
#10;
address_ina = 50;
address_inb = 51;
data_ina = 16'h193;
data_inb = 16'h5d7;
#10;
address_ina = 52;
address_inb = 53;
data_ina = 16'hfd89;
data_inb = 16'h294;
#10;
address_ina = 54;
address_inb = 55;
data_ina = 16'h577;
data_inb = 16'hfbc5;
#10;
address_ina = 56;
address_inb = 57;
data_ina = 16'hc9;
data_inb = 16'hfd6b;
#10;
address_ina = 58;
address_inb = 59;
data_ina = 16'h1f0;
data_inb = 16'h472;
#10;
address_ina = 60;
address_inb = 61;
data_ina = 16'h5c9;
data_inb = 16'h5d9;
#10;
address_ina = 62;
address_inb = 63;
data_ina = 16'hfcb0;
data_inb = 16'h3cf;
#10;
address_ina = 64;
address_inb = 65;
data_ina = 16'hfe61;
data_inb = 16'hfef8;
#10;
address_ina = 66;
address_inb = 67;
data_ina = 16'h176;
data_inb = 16'hfbff;
#10;
address_ina = 68;
address_inb = 69;
data_ina = 16'h1df;
data_inb = 16'h4b2;
#10;
address_ina = 70;
address_inb = 71;
data_ina = 16'hfacd;
data_inb = 16'h1e8;
#10;
address_ina = 72;
address_inb = 73;
data_ina = 16'h5d2;
data_inb = 16'h2d6;
#10;
address_ina = 74;
address_inb = 75;
data_ina = 16'h144;
data_inb = 16'hfcd8;
#10;
address_ina = 76;
address_inb = 77;
data_ina = 16'h8e;
data_inb = 16'hf9d4;
#10;
address_ina = 78;
address_inb = 79;
data_ina = 16'hfb7d;
data_inb = 16'hf9ed;
#10;
address_ina = 80;
address_inb = 81;
data_ina = 16'hfd10;
data_inb = 16'hfc67;
#10;
address_ina = 82;
address_inb = 83;
data_ina = 16'hfe64;
data_inb = 16'hffa2;
#10;
address_ina = 84;
address_inb = 85;
data_ina = 16'h52d;
data_inb = 16'hea;
#10;
address_ina = 86;
address_inb = 87;
data_ina = 16'h37c;
data_inb = 16'hfebe;
#10;
address_ina = 88;
address_inb = 89;
data_ina = 16'h36a;
data_inb = 16'hfd33;
#10;
address_ina = 90;
address_inb = 91;
data_ina = 16'h158;
data_inb = 16'h30;
#10;
address_ina = 92;
address_inb = 93;
data_ina = 16'h618;
data_inb = 16'hfbb3;
#10;
address_ina = 94;
address_inb = 95;
data_ina = 16'hfdd2;
data_inb = 16'hfd1d;
#10;
address_ina = 96;
address_inb = 97;
data_ina = 16'hfc9a;
data_inb = 16'hfdec;
#10;
address_ina = 98;
address_inb = 99;
data_ina = 16'hfdd4;
data_inb = 16'hfe21;
#10;
address_ina = 100;
address_inb = 101;
data_ina = 16'h643;
data_inb = 16'hfbc5;
#10;
address_ina = 102;
address_inb = 103;
data_ina = 16'hfce2;
data_inb = 16'h206;
#10;
address_ina = 104;
address_inb = 105;
data_ina = 16'hfe00;
data_inb = 16'h2db;
#10;
address_ina = 106;
address_inb = 107;
data_ina = 16'h58;
data_inb = 16'h2e6;
#10;
address_ina = 108;
address_inb = 109;
data_ina = 16'hfb7c;
data_inb = 16'hfd14;
#10;
address_ina = 110;
address_inb = 111;
data_ina = 16'h430;
data_inb = 16'hfe9b;
#10;
address_ina = 112;
address_inb = 113;
data_ina = 16'hfa5a;
data_inb = 16'h31e;
#10;
address_ina = 114;
address_inb = 115;
data_ina = 16'h599;
data_inb = 16'h5a5;
#10;
address_ina = 116;
address_inb = 117;
data_ina = 16'h30b;
data_inb = 16'hfa56;
#10;
address_ina = 118;
address_inb = 119;
data_ina = 16'h573;
data_inb = 16'hfc3e;
#10;
address_ina = 120;
address_inb = 121;
data_ina = 16'hff62;
data_inb = 16'hfc69;
#10;
address_ina = 122;
address_inb = 123;
data_ina = 16'hf99d;
data_inb = 16'h654;
#10;
address_ina = 124;
address_inb = 125;
data_ina = 16'h3a9;
data_inb = 16'h322;
#10;
address_ina = 126;
address_inb = 127;
data_ina = 16'hfd6a;
data_inb = 16'hfa7c;
#10;
address_ina = 128;
address_inb = 129;
data_ina = 16'hfcc3;
data_inb = 16'hfe7f;
#10;
address_ina = 130;
address_inb = 131;
data_ina = 16'h403;
data_inb = 16'hfbde;
#10;
address_ina = 132;
address_inb = 133;
data_ina = 16'hfa89;
data_inb = 16'hfe2e;
#10;
address_ina = 134;
address_inb = 135;
data_ina = 16'hfe2d;
data_inb = 16'hfb0c;
#10;
address_ina = 136;
address_inb = 137;
data_ina = 16'h21e;
data_inb = 16'h58d;
#10;
address_ina = 138;
address_inb = 139;
data_ina = 16'h18d;
data_inb = 16'hfae9;
#10;
address_ina = 140;
address_inb = 141;
data_ina = 16'h7;
data_inb = 16'hfef8;
#10;
address_ina = 142;
address_inb = 143;
data_ina = 16'hfe1d;
data_inb = 16'h30f;
#10;
address_ina = 144;
address_inb = 145;
data_ina = 16'h11b;
data_inb = 16'h486;
#10;
address_ina = 146;
address_inb = 147;
data_ina = 16'hfcb6;
data_inb = 16'h43;
#10;
address_ina = 148;
address_inb = 149;
data_ina = 16'hfb43;
data_inb = 16'h243;
#10;
address_ina = 150;
address_inb = 151;
data_ina = 16'h84;
data_inb = 16'h555;
#10;
address_ina = 152;
address_inb = 153;
data_ina = 16'h372;
data_inb = 16'h222;
#10;
address_ina = 154;
address_inb = 155;
data_ina = 16'hfcd6;
data_inb = 16'hfe8b;
#10;
address_ina = 156;
address_inb = 157;
data_ina = 16'h5ef;
data_inb = 16'hfe51;
#10;
address_ina = 158;
address_inb = 159;
data_ina = 16'hfc24;
data_inb = 16'h1e;
#10;
address_ina = 160;
address_inb = 161;
data_ina = 16'h60e;
data_inb = 16'hff;
#10;
address_ina = 162;
address_inb = 163;
data_ina = 16'hfe1d;
data_inb = 16'h480;
#10;
address_ina = 164;
address_inb = 165;
data_ina = 16'hfc19;
data_inb = 16'hfcb5;
#10;
address_ina = 166;
address_inb = 167;
data_ina = 16'h221;
data_inb = 16'h43f;
#10;
address_ina = 168;
address_inb = 169;
data_ina = 16'hfccf;
data_inb = 16'hfc47;
#10;
address_ina = 170;
address_inb = 171;
data_ina = 16'h1fe;
data_inb = 16'hf9ff;
#10;
address_ina = 172;
address_inb = 173;
data_ina = 16'hfe38;
data_inb = 16'h5da;
#10;
address_ina = 174;
address_inb = 175;
data_ina = 16'h132;
data_inb = 16'hfdac;
#10;
address_ina = 176;
address_inb = 177;
data_ina = 16'h673;
data_inb = 16'hf9ba;
#10;
address_ina = 178;
address_inb = 179;
data_ina = 16'hfd19;
data_inb = 16'hfe72;
#10;
address_ina = 180;
address_inb = 181;
data_ina = 16'hfec3;
data_inb = 16'hfde6;
#10;
address_ina = 182;
address_inb = 183;
data_ina = 16'hfcd6;
data_inb = 16'h390;
#10;
address_ina = 184;
address_inb = 185;
data_ina = 16'hfd26;
data_inb = 16'h372;
#10;
address_ina = 186;
address_inb = 187;
data_ina = 16'h50b;
data_inb = 16'h248;
#10;
address_ina = 188;
address_inb = 189;
data_ina = 16'h4f4;
data_inb = 16'h88;
#10;
address_ina = 190;
address_inb = 191;
data_ina = 16'h3ed;
data_inb = 16'h1b1;
#10;
address_ina = 192;
address_inb = 193;
data_ina = 16'h5b8;
data_inb = 16'h81;
#10;
address_ina = 194;
address_inb = 195;
data_ina = 16'hfc53;
data_inb = 16'h546;
#10;
address_ina = 196;
address_inb = 197;
data_ina = 16'h3c9;
data_inb = 16'h3e9;
#10;
address_ina = 198;
address_inb = 199;
data_ina = 16'hf994;
data_inb = 16'h4da;
#10;
address_ina = 200;
address_inb = 201;
data_ina = 16'hfa89;
data_inb = 16'hfe0f;
#10;
address_ina = 202;
address_inb = 203;
data_ina = 16'h4a5;
data_inb = 16'hfb53;
#10;
address_ina = 204;
address_inb = 205;
data_ina = 16'h1be;
data_inb = 16'hff81;
#10;
address_ina = 206;
address_inb = 207;
data_ina = 16'hfa35;
data_inb = 16'h314;
#10;
address_ina = 208;
address_inb = 209;
data_ina = 16'hfdec;
data_inb = 16'h343;
#10;
address_ina = 210;
address_inb = 211;
data_ina = 16'h552;
data_inb = 16'h25;
#10;
address_ina = 212;
address_inb = 213;
data_ina = 16'h51d;
data_inb = 16'hff40;
#10;
address_ina = 214;
address_inb = 215;
data_ina = 16'h551;
data_inb = 16'hfc2a;
#10;
address_ina = 216;
address_inb = 217;
data_ina = 16'h5d3;
data_inb = 16'h5be;
#10;
address_ina = 218;
address_inb = 219;
data_ina = 16'h50a;
data_inb = 16'hfa32;
#10;
address_ina = 220;
address_inb = 221;
data_ina = 16'hb3;
data_inb = 16'h158;
#10;
address_ina = 222;
address_inb = 223;
data_ina = 16'hfcc0;
data_inb = 16'hfb26;
#10;
address_ina = 224;
address_inb = 225;
data_ina = 16'h5a0;
data_inb = 16'hfbaf;
#10;
address_ina = 226;
address_inb = 227;
data_ina = 16'hfdeb;
data_inb = 16'hf9dc;
#10;
address_ina = 228;
address_inb = 229;
data_ina = 16'hfadd;
data_inb = 16'hff33;
#10;
address_ina = 230;
address_inb = 231;
data_ina = 16'hfcaa;
data_inb = 16'hff13;
#10;
address_ina = 232;
address_inb = 233;
data_ina = 16'h335;
data_inb = 16'h3e3;
#10;
address_ina = 234;
address_inb = 235;
data_ina = 16'hf9e4;
data_inb = 16'hfe1e;
#10;
address_ina = 236;
address_inb = 237;
data_ina = 16'h322;
data_inb = 16'h5d1;
#10;
address_ina = 238;
address_inb = 239;
data_ina = 16'h3f7;
data_inb = 16'hfb19;
#10;
address_ina = 240;
address_inb = 241;
data_ina = 16'hfd19;
data_inb = 16'hfc38;
#10;
address_ina = 242;
address_inb = 243;
data_ina = 16'h48c;
data_inb = 16'h45d;
#10;
address_ina = 244;
address_inb = 245;
data_ina = 16'hfb1a;
data_inb = 16'h4d6;
#10;
address_ina = 246;
address_inb = 247;
data_ina = 16'h101;
data_inb = 16'hfae1;
#10;
address_ina = 248;
address_inb = 249;
data_ina = 16'hfc18;
data_inb = 16'h369;
#10;
address_ina = 250;
address_inb = 251;
data_ina = 16'h1b0;
data_inb = 16'h185;
#10;
address_ina = 252;
address_inb = 253;
data_ina = 16'h28f;
data_inb = 16'hfae9;
#10;
address_ina = 254;
address_inb = 255;
data_ina = 16'hfbc0;
data_inb = 16'h2b4;
#10;
        wait(init_done);
        #30
        we = 0;
        // Start processing
         
		  #38000

        start = 0;



//        wait (wr_req);
//		  wait (!wr_req);
//		   rd_req = 1;
		  wait(done);
		  #20000
rd_req = 1;
        #70 
		  start = 1;
		 #80 
wait(rd_empty)
rd_req = 0;

$display("Finished the NTT test Number %d",test_num);
////Begin test number #41//////////////
rst = 1;

//#1000
start = 1;
mode = 1; //NTT 0 // INTT 1

// Reset for a few clock cycles

#1000

rst = 0;
test_num = test_num + 1;
#1000
we = 1;
address_ina = 0;
address_inb = 1;
data_ina = 16'h582;
data_inb = 16'hfa79;
#10;
address_ina = 2;
address_inb = 3;
data_ina = 16'hfd8d;
data_inb = 16'hfad4;
#10;
address_ina = 4;
address_inb = 5;
data_ina = 16'h1b8;
data_inb = 16'hff;
#10;
address_ina = 6;
address_inb = 7;
data_ina = 16'hfa3c;
data_inb = 16'h3d2;
#10;
address_ina = 8;
address_inb = 9;
data_ina = 16'hff83;
data_inb = 16'h460;
#10;
address_ina = 10;
address_inb = 11;
data_ina = 16'hfdb0;
data_inb = 16'h5a3;
#10;
address_ina = 12;
address_inb = 13;
data_ina = 16'h3b2;
data_inb = 16'hfdea;
#10;
address_ina = 14;
address_inb = 15;
data_ina = 16'hfb27;
data_inb = 16'h107;
#10;
address_ina = 16;
address_inb = 17;
data_ina = 16'hffbb;
data_inb = 16'h511;
#10;
address_ina = 18;
address_inb = 19;
data_ina = 16'h2b9;
data_inb = 16'hfcda;
#10;
address_ina = 20;
address_inb = 21;
data_ina = 16'hff35;
data_inb = 16'hfa9e;
#10;
address_ina = 22;
address_inb = 23;
data_ina = 16'hfc43;
data_inb = 16'hfd32;
#10;
address_ina = 24;
address_inb = 25;
data_ina = 16'h1d4;
data_inb = 16'hc6;
#10;
address_ina = 26;
address_inb = 27;
data_ina = 16'hfe27;
data_inb = 16'h557;
#10;
address_ina = 28;
address_inb = 29;
data_ina = 16'hfb2c;
data_inb = 16'h318;
#10;
address_ina = 30;
address_inb = 31;
data_ina = 16'h1f8;
data_inb = 16'hfe2b;
#10;
address_ina = 32;
address_inb = 33;
data_ina = 16'h633;
data_inb = 16'hfbcd;
#10;
address_ina = 34;
address_inb = 35;
data_ina = 16'hf9f8;
data_inb = 16'h41f;
#10;
address_ina = 36;
address_inb = 37;
data_ina = 16'hfe9d;
data_inb = 16'h35c;
#10;
address_ina = 38;
address_inb = 39;
data_ina = 16'h1c7;
data_inb = 16'h35f;
#10;
address_ina = 40;
address_inb = 41;
data_ina = 16'h637;
data_inb = 16'h57;
#10;
address_ina = 42;
address_inb = 43;
data_ina = 16'h313;
data_inb = 16'hfc2d;
#10;
address_ina = 44;
address_inb = 45;
data_ina = 16'ha2;
data_inb = 16'h65c;
#10;
address_ina = 46;
address_inb = 47;
data_ina = 16'h326;
data_inb = 16'hf9c0;
#10;
address_ina = 48;
address_inb = 49;
data_ina = 16'h4e4;
data_inb = 16'h4fc;
#10;
address_ina = 50;
address_inb = 51;
data_ina = 16'hfc01;
data_inb = 16'hfaa5;
#10;
address_ina = 52;
address_inb = 53;
data_ina = 16'h62d;
data_inb = 16'hfda0;
#10;
address_ina = 54;
address_inb = 55;
data_ina = 16'h662;
data_inb = 16'h44d;
#10;
address_ina = 56;
address_inb = 57;
data_ina = 16'hf9d0;
data_inb = 16'hdb;
#10;
address_ina = 58;
address_inb = 59;
data_ina = 16'hf984;
data_inb = 16'h37f;
#10;
address_ina = 60;
address_inb = 61;
data_ina = 16'hf9cf;
data_inb = 16'h2b4;
#10;
address_ina = 62;
address_inb = 63;
data_ina = 16'hfd59;
data_inb = 16'hfe0f;
#10;
address_ina = 64;
address_inb = 65;
data_ina = 16'h62b;
data_inb = 16'h4ee;
#10;
address_ina = 66;
address_inb = 67;
data_ina = 16'hfc5e;
data_inb = 16'h504;
#10;
address_ina = 68;
address_inb = 69;
data_ina = 16'hffab;
data_inb = 16'hff08;
#10;
address_ina = 70;
address_inb = 71;
data_ina = 16'h23c;
data_inb = 16'hfc1f;
#10;
address_ina = 72;
address_inb = 73;
data_ina = 16'hfe6c;
data_inb = 16'h5dc;
#10;
address_ina = 74;
address_inb = 75;
data_ina = 16'hfea1;
data_inb = 16'h5d3;
#10;
address_ina = 76;
address_inb = 77;
data_ina = 16'hc8;
data_inb = 16'hf9df;
#10;
address_ina = 78;
address_inb = 79;
data_ina = 16'h40d;
data_inb = 16'h512;
#10;
address_ina = 80;
address_inb = 81;
data_ina = 16'h616;
data_inb = 16'hfe57;
#10;
address_ina = 82;
address_inb = 83;
data_ina = 16'hfc44;
data_inb = 16'h95;
#10;
address_ina = 84;
address_inb = 85;
data_ina = 16'hfc90;
data_inb = 16'hfb66;
#10;
address_ina = 86;
address_inb = 87;
data_ina = 16'h35d;
data_inb = 16'h45b;
#10;
address_ina = 88;
address_inb = 89;
data_ina = 16'hfdac;
data_inb = 16'h2bb;
#10;
address_ina = 90;
address_inb = 91;
data_ina = 16'h90;
data_inb = 16'h138;
#10;
address_ina = 92;
address_inb = 93;
data_ina = 16'hfbc8;
data_inb = 16'h5c0;
#10;
address_ina = 94;
address_inb = 95;
data_ina = 16'h58;
data_inb = 16'hfe0b;
#10;
address_ina = 96;
address_inb = 97;
data_ina = 16'hfe8b;
data_inb = 16'hffe0;
#10;
address_ina = 98;
address_inb = 99;
data_ina = 16'hffd8;
data_inb = 16'hfdaf;
#10;
address_ina = 100;
address_inb = 101;
data_ina = 16'h5e2;
data_inb = 16'hfd95;
#10;
address_ina = 102;
address_inb = 103;
data_ina = 16'hfc71;
data_inb = 16'hfdb9;
#10;
address_ina = 104;
address_inb = 105;
data_ina = 16'h5a7;
data_inb = 16'hffea;
#10;
address_ina = 106;
address_inb = 107;
data_ina = 16'h3e7;
data_inb = 16'h2a8;
#10;
address_ina = 108;
address_inb = 109;
data_ina = 16'h51c;
data_inb = 16'hfc74;
#10;
address_ina = 110;
address_inb = 111;
data_ina = 16'hfcc7;
data_inb = 16'h4dd;
#10;
address_ina = 112;
address_inb = 113;
data_ina = 16'h5ad;
data_inb = 16'hfc3c;
#10;
address_ina = 114;
address_inb = 115;
data_ina = 16'hfd9d;
data_inb = 16'h52c;
#10;
address_ina = 116;
address_inb = 117;
data_ina = 16'h16b;
data_inb = 16'hffcb;
#10;
address_ina = 118;
address_inb = 119;
data_ina = 16'hfcfc;
data_inb = 16'hfb6e;
#10;
address_ina = 120;
address_inb = 121;
data_ina = 16'hfd55;
data_inb = 16'hfa58;
#10;
address_ina = 122;
address_inb = 123;
data_ina = 16'hfb29;
data_inb = 16'h35a;
#10;
address_ina = 124;
address_inb = 125;
data_ina = 16'h474;
data_inb = 16'h2e8;
#10;
address_ina = 126;
address_inb = 127;
data_ina = 16'h298;
data_inb = 16'hfcc8;
#10;
address_ina = 128;
address_inb = 129;
data_ina = 16'hfc71;
data_inb = 16'hfd66;
#10;
address_ina = 130;
address_inb = 131;
data_ina = 16'h4e3;
data_inb = 16'hfacb;
#10;
address_ina = 132;
address_inb = 133;
data_ina = 16'hf9ae;
data_inb = 16'h5b2;
#10;
address_ina = 134;
address_inb = 135;
data_ina = 16'h49d;
data_inb = 16'h457;
#10;
address_ina = 136;
address_inb = 137;
data_ina = 16'hffeb;
data_inb = 16'h328;
#10;
address_ina = 138;
address_inb = 139;
data_ina = 16'h3ec;
data_inb = 16'hfd4e;
#10;
address_ina = 140;
address_inb = 141;
data_ina = 16'h418;
data_inb = 16'hfc63;
#10;
address_ina = 142;
address_inb = 143;
data_ina = 16'h1a8;
data_inb = 16'h44a;
#10;
address_ina = 144;
address_inb = 145;
data_ina = 16'hff95;
data_inb = 16'hfc62;
#10;
address_ina = 146;
address_inb = 147;
data_ina = 16'h42f;
data_inb = 16'h624;
#10;
address_ina = 148;
address_inb = 149;
data_ina = 16'hfdfe;
data_inb = 16'h388;
#10;
address_ina = 150;
address_inb = 151;
data_ina = 16'hfc7d;
data_inb = 16'h64e;
#10;
address_ina = 152;
address_inb = 153;
data_ina = 16'hfe3a;
data_inb = 16'h1ce;
#10;
address_ina = 154;
address_inb = 155;
data_ina = 16'hfe94;
data_inb = 16'hfc34;
#10;
address_ina = 156;
address_inb = 157;
data_ina = 16'hff07;
data_inb = 16'hfcb1;
#10;
address_ina = 158;
address_inb = 159;
data_ina = 16'hfc46;
data_inb = 16'h157;
#10;
address_ina = 160;
address_inb = 161;
data_ina = 16'h1e6;
data_inb = 16'hfdb3;
#10;
address_ina = 162;
address_inb = 163;
data_ina = 16'hfda7;
data_inb = 16'hfb81;
#10;
address_ina = 164;
address_inb = 165;
data_ina = 16'hf9d4;
data_inb = 16'hfb88;
#10;
address_ina = 166;
address_inb = 167;
data_ina = 16'hfe79;
data_inb = 16'h488;
#10;
address_ina = 168;
address_inb = 169;
data_ina = 16'hfebc;
data_inb = 16'hfeb1;
#10;
address_ina = 170;
address_inb = 171;
data_ina = 16'hfbe4;
data_inb = 16'hfe78;
#10;
address_ina = 172;
address_inb = 173;
data_ina = 16'h67d;
data_inb = 16'h3ed;
#10;
address_ina = 174;
address_inb = 175;
data_ina = 16'h1c0;
data_inb = 16'hffe5;
#10;
address_ina = 176;
address_inb = 177;
data_ina = 16'hfebd;
data_inb = 16'h3ba;
#10;
address_ina = 178;
address_inb = 179;
data_ina = 16'hfc96;
data_inb = 16'hff5e;
#10;
address_ina = 180;
address_inb = 181;
data_ina = 16'hfcad;
data_inb = 16'hfffe;
#10;
address_ina = 182;
address_inb = 183;
data_ina = 16'hfb4c;
data_inb = 16'h644;
#10;
address_ina = 184;
address_inb = 185;
data_ina = 16'hf9d3;
data_inb = 16'hff49;
#10;
address_ina = 186;
address_inb = 187;
data_ina = 16'h3dc;
data_inb = 16'hfae8;
#10;
address_ina = 188;
address_inb = 189;
data_ina = 16'h4d5;
data_inb = 16'hff88;
#10;
address_ina = 190;
address_inb = 191;
data_ina = 16'h37a;
data_inb = 16'h3f2;
#10;
address_ina = 192;
address_inb = 193;
data_ina = 16'h104;
data_inb = 16'h5f1;
#10;
address_ina = 194;
address_inb = 195;
data_ina = 16'hfa87;
data_inb = 16'hff6c;
#10;
address_ina = 196;
address_inb = 197;
data_ina = 16'h429;
data_inb = 16'h1a1;
#10;
address_ina = 198;
address_inb = 199;
data_ina = 16'hffe5;
data_inb = 16'hfcae;
#10;
address_ina = 200;
address_inb = 201;
data_ina = 16'hfd88;
data_inb = 16'h3ad;
#10;
address_ina = 202;
address_inb = 203;
data_ina = 16'hfd13;
data_inb = 16'hff97;
#10;
address_ina = 204;
address_inb = 205;
data_ina = 16'hfec5;
data_inb = 16'hc3;
#10;
address_ina = 206;
address_inb = 207;
data_ina = 16'h42c;
data_inb = 16'hfb68;
#10;
address_ina = 208;
address_inb = 209;
data_ina = 16'h34;
data_inb = 16'h274;
#10;
address_ina = 210;
address_inb = 211;
data_ina = 16'hfca0;
data_inb = 16'h641;
#10;
address_ina = 212;
address_inb = 213;
data_ina = 16'h4c9;
data_inb = 16'h431;
#10;
address_ina = 214;
address_inb = 215;
data_ina = 16'h50b;
data_inb = 16'h669;
#10;
address_ina = 216;
address_inb = 217;
data_ina = 16'hfdaf;
data_inb = 16'h3ec;
#10;
address_ina = 218;
address_inb = 219;
data_ina = 16'h2a3;
data_inb = 16'hfe59;
#10;
address_ina = 220;
address_inb = 221;
data_ina = 16'h332;
data_inb = 16'h11c;
#10;
address_ina = 222;
address_inb = 223;
data_ina = 16'hfa04;
data_inb = 16'h568;
#10;
address_ina = 224;
address_inb = 225;
data_ina = 16'hf9b0;
data_inb = 16'hfd29;
#10;
address_ina = 226;
address_inb = 227;
data_ina = 16'h438;
data_inb = 16'hfee8;
#10;
address_ina = 228;
address_inb = 229;
data_ina = 16'h635;
data_inb = 16'h17d;
#10;
address_ina = 230;
address_inb = 231;
data_ina = 16'hfa0c;
data_inb = 16'h3bc;
#10;
address_ina = 232;
address_inb = 233;
data_ina = 16'hffa7;
data_inb = 16'h49f;
#10;
address_ina = 234;
address_inb = 235;
data_ina = 16'hfacc;
data_inb = 16'hfd00;
#10;
address_ina = 236;
address_inb = 237;
data_ina = 16'h40;
data_inb = 16'hf99c;
#10;
address_ina = 238;
address_inb = 239;
data_ina = 16'hfdec;
data_inb = 16'ha9;
#10;
address_ina = 240;
address_inb = 241;
data_ina = 16'hff07;
data_inb = 16'hffe6;
#10;
address_ina = 242;
address_inb = 243;
data_ina = 16'h613;
data_inb = 16'hfe14;
#10;
address_ina = 244;
address_inb = 245;
data_ina = 16'hfa42;
data_inb = 16'h13d;
#10;
address_ina = 246;
address_inb = 247;
data_ina = 16'h4a;
data_inb = 16'h309;
#10;
address_ina = 248;
address_inb = 249;
data_ina = 16'hf9a4;
data_inb = 16'hfdbb;
#10;
address_ina = 250;
address_inb = 251;
data_ina = 16'hb5;
data_inb = 16'h24c;
#10;
address_ina = 252;
address_inb = 253;
data_ina = 16'h252;
data_inb = 16'h449;
#10;
address_ina = 254;
address_inb = 255;
data_ina = 16'h3d3;
data_inb = 16'hfcc2;
#10;
        wait(init_done);
        #30
        we = 0;
        // Start processing
         
		  #38000

        start = 0;



//        wait (wr_req);
//		  wait (!wr_req);
//		   rd_req = 1;
		  wait(done);
		  #20000
rd_req = 1;
        #70 
		  start = 1;
		 #80 
wait(rd_empty)
rd_req = 0;

$display("Finished the NTT test Number %d",test_num);
////Begin test number #42//////////////
rst = 1;

//#1000
start = 1;
mode = 1; //NTT 0 // INTT 1

// Reset for a few clock cycles

#1000

rst = 0;
test_num = test_num + 1;
#1000
we = 1;
address_ina = 0;
address_inb = 1;
data_ina = 16'hff21;
data_inb = 16'hfa22;
#10;
address_ina = 2;
address_inb = 3;
data_ina = 16'h457;
data_inb = 16'hfecc;
#10;
address_ina = 4;
address_inb = 5;
data_ina = 16'hff3e;
data_inb = 16'hf9ab;
#10;
address_ina = 6;
address_inb = 7;
data_ina = 16'h2c9;
data_inb = 16'hfca2;
#10;
address_ina = 8;
address_inb = 9;
data_ina = 16'hfa45;
data_inb = 16'hfa84;
#10;
address_ina = 10;
address_inb = 11;
data_ina = 16'hfd99;
data_inb = 16'h4ca;
#10;
address_ina = 12;
address_inb = 13;
data_ina = 16'h364;
data_inb = 16'hfb9e;
#10;
address_ina = 14;
address_inb = 15;
data_ina = 16'h4b3;
data_inb = 16'hff77;
#10;
address_ina = 16;
address_inb = 17;
data_ina = 16'h9f;
data_inb = 16'hdc;
#10;
address_ina = 18;
address_inb = 19;
data_ina = 16'hfe5f;
data_inb = 16'hff51;
#10;
address_ina = 20;
address_inb = 21;
data_ina = 16'hfb5e;
data_inb = 16'hfac2;
#10;
address_ina = 22;
address_inb = 23;
data_ina = 16'hff43;
data_inb = 16'h596;
#10;
address_ina = 24;
address_inb = 25;
data_ina = 16'hff94;
data_inb = 16'hfa43;
#10;
address_ina = 26;
address_inb = 27;
data_ina = 16'h14e;
data_inb = 16'hffe2;
#10;
address_ina = 28;
address_inb = 29;
data_ina = 16'hfc8f;
data_inb = 16'h33c;
#10;
address_ina = 30;
address_inb = 31;
data_ina = 16'hfb1f;
data_inb = 16'h12c;
#10;
address_ina = 32;
address_inb = 33;
data_ina = 16'hfdec;
data_inb = 16'hfd50;
#10;
address_ina = 34;
address_inb = 35;
data_ina = 16'hf9b8;
data_inb = 16'h5bc;
#10;
address_ina = 36;
address_inb = 37;
data_ina = 16'hff19;
data_inb = 16'h403;
#10;
address_ina = 38;
address_inb = 39;
data_ina = 16'hfa7f;
data_inb = 16'hff6d;
#10;
address_ina = 40;
address_inb = 41;
data_ina = 16'h53d;
data_inb = 16'hfa1b;
#10;
address_ina = 42;
address_inb = 43;
data_ina = 16'h37;
data_inb = 16'hfa9c;
#10;
address_ina = 44;
address_inb = 45;
data_ina = 16'hfa32;
data_inb = 16'hfe0c;
#10;
address_ina = 46;
address_inb = 47;
data_ina = 16'hfb24;
data_inb = 16'h223;
#10;
address_ina = 48;
address_inb = 49;
data_ina = 16'hfcc0;
data_inb = 16'hffb1;
#10;
address_ina = 50;
address_inb = 51;
data_ina = 16'h48e;
data_inb = 16'h66f;
#10;
address_ina = 52;
address_inb = 53;
data_ina = 16'hfca5;
data_inb = 16'h1a4;
#10;
address_ina = 54;
address_inb = 55;
data_ina = 16'hfd5a;
data_inb = 16'h4d3;
#10;
address_ina = 56;
address_inb = 57;
data_ina = 16'h1d9;
data_inb = 16'h4e6;
#10;
address_ina = 58;
address_inb = 59;
data_ina = 16'hfc6b;
data_inb = 16'hfcb2;
#10;
address_ina = 60;
address_inb = 61;
data_ina = 16'hfdde;
data_inb = 16'hfdd6;
#10;
address_ina = 62;
address_inb = 63;
data_ina = 16'hfcb2;
data_inb = 16'h447;
#10;
address_ina = 64;
address_inb = 65;
data_ina = 16'h350;
data_inb = 16'hfcf4;
#10;
address_ina = 66;
address_inb = 67;
data_ina = 16'hf992;
data_inb = 16'h636;
#10;
address_ina = 68;
address_inb = 69;
data_ina = 16'h32f;
data_inb = 16'hfdb9;
#10;
address_ina = 70;
address_inb = 71;
data_ina = 16'h497;
data_inb = 16'h256;
#10;
address_ina = 72;
address_inb = 73;
data_ina = 16'hfdbe;
data_inb = 16'hfaa5;
#10;
address_ina = 74;
address_inb = 75;
data_ina = 16'hfaa5;
data_inb = 16'hfa40;
#10;
address_ina = 76;
address_inb = 77;
data_ina = 16'h13d;
data_inb = 16'h3e2;
#10;
address_ina = 78;
address_inb = 79;
data_ina = 16'hfdf3;
data_inb = 16'hfc0d;
#10;
address_ina = 80;
address_inb = 81;
data_ina = 16'h5c8;
data_inb = 16'hfc46;
#10;
address_ina = 82;
address_inb = 83;
data_ina = 16'hfa23;
data_inb = 16'h62a;
#10;
address_ina = 84;
address_inb = 85;
data_ina = 16'h3d6;
data_inb = 16'h272;
#10;
address_ina = 86;
address_inb = 87;
data_ina = 16'hfba0;
data_inb = 16'h58b;
#10;
address_ina = 88;
address_inb = 89;
data_ina = 16'hfd23;
data_inb = 16'h63e;
#10;
address_ina = 90;
address_inb = 91;
data_ina = 16'h69;
data_inb = 16'h521;
#10;
address_ina = 92;
address_inb = 93;
data_ina = 16'hbd;
data_inb = 16'hfcdd;
#10;
address_ina = 94;
address_inb = 95;
data_ina = 16'h524;
data_inb = 16'hfb5f;
#10;
address_ina = 96;
address_inb = 97;
data_ina = 16'hfbe0;
data_inb = 16'h5dd;
#10;
address_ina = 98;
address_inb = 99;
data_ina = 16'hfee2;
data_inb = 16'h2f6;
#10;
address_ina = 100;
address_inb = 101;
data_ina = 16'h181;
data_inb = 16'h611;
#10;
address_ina = 102;
address_inb = 103;
data_ina = 16'hff4b;
data_inb = 16'h291;
#10;
address_ina = 104;
address_inb = 105;
data_ina = 16'hf9d9;
data_inb = 16'hfad3;
#10;
address_ina = 106;
address_inb = 107;
data_ina = 16'hfda0;
data_inb = 16'h11;
#10;
address_ina = 108;
address_inb = 109;
data_ina = 16'hff67;
data_inb = 16'hfb80;
#10;
address_ina = 110;
address_inb = 111;
data_ina = 16'h505;
data_inb = 16'h597;
#10;
address_ina = 112;
address_inb = 113;
data_ina = 16'hffe5;
data_inb = 16'hfcb4;
#10;
address_ina = 114;
address_inb = 115;
data_ina = 16'h104;
data_inb = 16'h4c9;
#10;
address_ina = 116;
address_inb = 117;
data_ina = 16'h233;
data_inb = 16'hfccc;
#10;
address_ina = 118;
address_inb = 119;
data_ina = 16'h98;
data_inb = 16'hfab6;
#10;
address_ina = 120;
address_inb = 121;
data_ina = 16'hfe78;
data_inb = 16'h61f;
#10;
address_ina = 122;
address_inb = 123;
data_ina = 16'h182;
data_inb = 16'h1a;
#10;
address_ina = 124;
address_inb = 125;
data_ina = 16'h436;
data_inb = 16'h1b;
#10;
address_ina = 126;
address_inb = 127;
data_ina = 16'h5ce;
data_inb = 16'h498;
#10;
address_ina = 128;
address_inb = 129;
data_ina = 16'h71;
data_inb = 16'hfe4d;
#10;
address_ina = 130;
address_inb = 131;
data_ina = 16'h5a8;
data_inb = 16'h580;
#10;
address_ina = 132;
address_inb = 133;
data_ina = 16'h5bc;
data_inb = 16'h5ca;
#10;
address_ina = 134;
address_inb = 135;
data_ina = 16'hfe17;
data_inb = 16'hfdd0;
#10;
address_ina = 136;
address_inb = 137;
data_ina = 16'h385;
data_inb = 16'hfb32;
#10;
address_ina = 138;
address_inb = 139;
data_ina = 16'hfe63;
data_inb = 16'hf9e8;
#10;
address_ina = 140;
address_inb = 141;
data_ina = 16'h42e;
data_inb = 16'h458;
#10;
address_ina = 142;
address_inb = 143;
data_ina = 16'hff02;
data_inb = 16'hf9a0;
#10;
address_ina = 144;
address_inb = 145;
data_ina = 16'hffb2;
data_inb = 16'hfe18;
#10;
address_ina = 146;
address_inb = 147;
data_ina = 16'hfd9a;
data_inb = 16'h38d;
#10;
address_ina = 148;
address_inb = 149;
data_ina = 16'hfaed;
data_inb = 16'hfb01;
#10;
address_ina = 150;
address_inb = 151;
data_ina = 16'hf9da;
data_inb = 16'h322;
#10;
address_ina = 152;
address_inb = 153;
data_ina = 16'hf9f1;
data_inb = 16'hffd3;
#10;
address_ina = 154;
address_inb = 155;
data_ina = 16'h47c;
data_inb = 16'hfa2b;
#10;
address_ina = 156;
address_inb = 157;
data_ina = 16'h69;
data_inb = 16'h4ee;
#10;
address_ina = 158;
address_inb = 159;
data_ina = 16'hfd7f;
data_inb = 16'hfb14;
#10;
address_ina = 160;
address_inb = 161;
data_ina = 16'hff2e;
data_inb = 16'hfcb6;
#10;
address_ina = 162;
address_inb = 163;
data_ina = 16'hfaf1;
data_inb = 16'hffd8;
#10;
address_ina = 164;
address_inb = 165;
data_ina = 16'hfdeb;
data_inb = 16'hfd29;
#10;
address_ina = 166;
address_inb = 167;
data_ina = 16'h418;
data_inb = 16'ha5;
#10;
address_ina = 168;
address_inb = 169;
data_ina = 16'hfa12;
data_inb = 16'hfbdc;
#10;
address_ina = 170;
address_inb = 171;
data_ina = 16'h4a9;
data_inb = 16'hff9e;
#10;
address_ina = 172;
address_inb = 173;
data_ina = 16'hfdd1;
data_inb = 16'hfa04;
#10;
address_ina = 174;
address_inb = 175;
data_ina = 16'h47a;
data_inb = 16'hff27;
#10;
address_ina = 176;
address_inb = 177;
data_ina = 16'h5f6;
data_inb = 16'h3a;
#10;
address_ina = 178;
address_inb = 179;
data_ina = 16'h20d;
data_inb = 16'hfd8b;
#10;
address_ina = 180;
address_inb = 181;
data_ina = 16'h4c0;
data_inb = 16'hfc7c;
#10;
address_ina = 182;
address_inb = 183;
data_ina = 16'hfd5d;
data_inb = 16'hfa92;
#10;
address_ina = 184;
address_inb = 185;
data_ina = 16'hfb59;
data_inb = 16'hfdf3;
#10;
address_ina = 186;
address_inb = 187;
data_ina = 16'h4f8;
data_inb = 16'hfe9c;
#10;
address_ina = 188;
address_inb = 189;
data_ina = 16'hfbc8;
data_inb = 16'h522;
#10;
address_ina = 190;
address_inb = 191;
data_ina = 16'hfbbc;
data_inb = 16'hff76;
#10;
address_ina = 192;
address_inb = 193;
data_ina = 16'h3d1;
data_inb = 16'h497;
#10;
address_ina = 194;
address_inb = 195;
data_ina = 16'ha3;
data_inb = 16'h17;
#10;
address_ina = 196;
address_inb = 197;
data_ina = 16'h5de;
data_inb = 16'h107;
#10;
address_ina = 198;
address_inb = 199;
data_ina = 16'hfac8;
data_inb = 16'h46c;
#10;
address_ina = 200;
address_inb = 201;
data_ina = 16'hd2;
data_inb = 16'hff1a;
#10;
address_ina = 202;
address_inb = 203;
data_ina = 16'hff0c;
data_inb = 16'hfaa2;
#10;
address_ina = 204;
address_inb = 205;
data_ina = 16'hfef1;
data_inb = 16'he8;
#10;
address_ina = 206;
address_inb = 207;
data_ina = 16'hffba;
data_inb = 16'hc8;
#10;
address_ina = 208;
address_inb = 209;
data_ina = 16'hfedd;
data_inb = 16'h158;
#10;
address_ina = 210;
address_inb = 211;
data_ina = 16'h63c;
data_inb = 16'hd6;
#10;
address_ina = 212;
address_inb = 213;
data_ina = 16'h4ae;
data_inb = 16'hfd17;
#10;
address_ina = 214;
address_inb = 215;
data_ina = 16'h137;
data_inb = 16'hf9b4;
#10;
address_ina = 216;
address_inb = 217;
data_ina = 16'hfda5;
data_inb = 16'hf99c;
#10;
address_ina = 218;
address_inb = 219;
data_ina = 16'h7c;
data_inb = 16'h62f;
#10;
address_ina = 220;
address_inb = 221;
data_ina = 16'h1e3;
data_inb = 16'hf99a;
#10;
address_ina = 222;
address_inb = 223;
data_ina = 16'h178;
data_inb = 16'hfd83;
#10;
address_ina = 224;
address_inb = 225;
data_ina = 16'he9;
data_inb = 16'h627;
#10;
address_ina = 226;
address_inb = 227;
data_ina = 16'hf9db;
data_inb = 16'ha8;
#10;
address_ina = 228;
address_inb = 229;
data_ina = 16'hfd0e;
data_inb = 16'h24a;
#10;
address_ina = 230;
address_inb = 231;
data_ina = 16'hfe5c;
data_inb = 16'h2e2;
#10;
address_ina = 232;
address_inb = 233;
data_ina = 16'hfb28;
data_inb = 16'h55f;
#10;
address_ina = 234;
address_inb = 235;
data_ina = 16'h23b;
data_inb = 16'hf980;
#10;
address_ina = 236;
address_inb = 237;
data_ina = 16'hfb33;
data_inb = 16'hfe36;
#10;
address_ina = 238;
address_inb = 239;
data_ina = 16'h154;
data_inb = 16'h66b;
#10;
address_ina = 240;
address_inb = 241;
data_ina = 16'hff78;
data_inb = 16'h2f;
#10;
address_ina = 242;
address_inb = 243;
data_ina = 16'h60a;
data_inb = 16'hfd43;
#10;
address_ina = 244;
address_inb = 245;
data_ina = 16'h7c;
data_inb = 16'h4ed;
#10;
address_ina = 246;
address_inb = 247;
data_ina = 16'hff7c;
data_inb = 16'h74;
#10;
address_ina = 248;
address_inb = 249;
data_ina = 16'h1fd;
data_inb = 16'hfab9;
#10;
address_ina = 250;
address_inb = 251;
data_ina = 16'hfb9a;
data_inb = 16'hff50;
#10;
address_ina = 252;
address_inb = 253;
data_ina = 16'h610;
data_inb = 16'hfa1a;
#10;
address_ina = 254;
address_inb = 255;
data_ina = 16'hff0c;
data_inb = 16'h494;
#10;
        wait(init_done);
        #30
        we = 0;
        // Start processing
         
		  #38000

        start = 0;



//        wait (wr_req);
//		  wait (!wr_req);
//		   rd_req = 1;
		  wait(done);
		  #20000
rd_req = 1;
        #70 
		  start = 1;
		 #80 
wait(rd_empty)
rd_req = 0;

$display("Finished the NTT test Number %d",test_num);
////Begin test number #43//////////////
rst = 1;

//#1000
start = 1;
mode = 0; //NTT 0 // INTT 1

// Reset for a few clock cycles

#1000

rst = 0;
test_num = test_num + 1;
#1000
we = 1;
address_ina = 0;
address_inb = 1;
data_ina = 16'hc85;
data_inb = 16'h4b6;
#10;
address_ina = 2;
address_inb = 3;
data_ina = 16'h2e2;
data_inb = 16'h618;
#10;
address_ina = 4;
address_inb = 5;
data_ina = 16'ha39;
data_inb = 16'h319;
#10;
address_ina = 6;
address_inb = 7;
data_ina = 16'h5ee;
data_inb = 16'h555;
#10;
address_ina = 8;
address_inb = 9;
data_ina = 16'h6f6;
data_inb = 16'h212;
#10;
address_ina = 10;
address_inb = 11;
data_ina = 16'h10b;
data_inb = 16'h8f;
#10;
address_ina = 12;
address_inb = 13;
data_ina = 16'h10e;
data_inb = 16'h6e9;
#10;
address_ina = 14;
address_inb = 15;
data_ina = 16'h3b9;
data_inb = 16'h1b0;
#10;
address_ina = 16;
address_inb = 17;
data_ina = 16'h180;
data_inb = 16'h754;
#10;
address_ina = 18;
address_inb = 19;
data_ina = 16'h294;
data_inb = 16'h14c;
#10;
address_ina = 20;
address_inb = 21;
data_ina = 16'hae9;
data_inb = 16'hb47;
#10;
address_ina = 22;
address_inb = 23;
data_ina = 16'hb26;
data_inb = 16'h398;
#10;
address_ina = 24;
address_inb = 25;
data_ina = 16'h1c4;
data_inb = 16'ha91;
#10;
address_ina = 26;
address_inb = 27;
data_ina = 16'h9c7;
data_inb = 16'h1c1;
#10;
address_ina = 28;
address_inb = 29;
data_ina = 16'h1fb;
data_inb = 16'h15c;
#10;
address_ina = 30;
address_inb = 31;
data_ina = 16'hbe6;
data_inb = 16'h882;
#10;
address_ina = 32;
address_inb = 33;
data_ina = 16'h4e7;
data_inb = 16'h542;
#10;
address_ina = 34;
address_inb = 35;
data_ina = 16'h767;
data_inb = 16'h80d;
#10;
address_ina = 36;
address_inb = 37;
data_ina = 16'h59d;
data_inb = 16'h875;
#10;
address_ina = 38;
address_inb = 39;
data_ina = 16'ha26;
data_inb = 16'h5b4;
#10;
address_ina = 40;
address_inb = 41;
data_ina = 16'hc21;
data_inb = 16'h3d3;
#10;
address_ina = 42;
address_inb = 43;
data_ina = 16'h58;
data_inb = 16'h4c6;
#10;
address_ina = 44;
address_inb = 45;
data_ina = 16'h1fe;
data_inb = 16'hbdc;
#10;
address_ina = 46;
address_inb = 47;
data_ina = 16'h263;
data_inb = 16'h7fd;
#10;
address_ina = 48;
address_inb = 49;
data_ina = 16'h72a;
data_inb = 16'h75a;
#10;
address_ina = 50;
address_inb = 51;
data_ina = 16'hb92;
data_inb = 16'h720;
#10;
address_ina = 52;
address_inb = 53;
data_ina = 16'h21;
data_inb = 16'h24;
#10;
address_ina = 54;
address_inb = 55;
data_ina = 16'h29a;
data_inb = 16'hb3a;
#10;
address_ina = 56;
address_inb = 57;
data_ina = 16'h259;
data_inb = 16'h273;
#10;
address_ina = 58;
address_inb = 59;
data_ina = 16'h5d1;
data_inb = 16'h1d4;
#10;
address_ina = 60;
address_inb = 61;
data_ina = 16'hc99;
data_inb = 16'h3e3;
#10;
address_ina = 62;
address_inb = 63;
data_ina = 16'h824;
data_inb = 16'h444;
#10;
address_ina = 64;
address_inb = 65;
data_ina = 16'h97c;
data_inb = 16'h9a0;
#10;
address_ina = 66;
address_inb = 67;
data_ina = 16'h7ac;
data_inb = 16'h969;
#10;
address_ina = 68;
address_inb = 69;
data_ina = 16'hca3;
data_inb = 16'h2a;
#10;
address_ina = 70;
address_inb = 71;
data_ina = 16'haa8;
data_inb = 16'hcea;
#10;
address_ina = 72;
address_inb = 73;
data_ina = 16'h586;
data_inb = 16'h37e;
#10;
address_ina = 74;
address_inb = 75;
data_ina = 16'ha;
data_inb = 16'h68a;
#10;
address_ina = 76;
address_inb = 77;
data_ina = 16'h848;
data_inb = 16'h8bd;
#10;
address_ina = 78;
address_inb = 79;
data_ina = 16'h444;
data_inb = 16'h329;
#10;
address_ina = 80;
address_inb = 81;
data_ina = 16'h2b4;
data_inb = 16'h5f1;
#10;
address_ina = 82;
address_inb = 83;
data_ina = 16'hcc3;
data_inb = 16'h771;
#10;
address_ina = 84;
address_inb = 85;
data_ina = 16'h986;
data_inb = 16'h256;
#10;
address_ina = 86;
address_inb = 87;
data_ina = 16'h4fa;
data_inb = 16'h458;
#10;
address_ina = 88;
address_inb = 89;
data_ina = 16'hb09;
data_inb = 16'ha26;
#10;
address_ina = 90;
address_inb = 91;
data_ina = 16'hbc9;
data_inb = 16'h2f2;
#10;
address_ina = 92;
address_inb = 93;
data_ina = 16'h94f;
data_inb = 16'h800;
#10;
address_ina = 94;
address_inb = 95;
data_ina = 16'h986;
data_inb = 16'h410;
#10;
address_ina = 96;
address_inb = 97;
data_ina = 16'h12b;
data_inb = 16'h50b;
#10;
address_ina = 98;
address_inb = 99;
data_ina = 16'hbe3;
data_inb = 16'ha0c;
#10;
address_ina = 100;
address_inb = 101;
data_ina = 16'h4e0;
data_inb = 16'h925;
#10;
address_ina = 102;
address_inb = 103;
data_ina = 16'hb26;
data_inb = 16'hcca;
#10;
address_ina = 104;
address_inb = 105;
data_ina = 16'h4b6;
data_inb = 16'h91e;
#10;
address_ina = 106;
address_inb = 107;
data_ina = 16'h354;
data_inb = 16'ha53;
#10;
address_ina = 108;
address_inb = 109;
data_ina = 16'h9ad;
data_inb = 16'hb40;
#10;
address_ina = 110;
address_inb = 111;
data_ina = 16'h270;
data_inb = 16'hc03;
#10;
address_ina = 112;
address_inb = 113;
data_ina = 16'h67d;
data_inb = 16'h40a;
#10;
address_ina = 114;
address_inb = 115;
data_ina = 16'h7dc;
data_inb = 16'hcea;
#10;
address_ina = 116;
address_inb = 117;
data_ina = 16'h1c1;
data_inb = 16'h41;
#10;
address_ina = 118;
address_inb = 119;
data_ina = 16'h6c5;
data_inb = 16'h309;
#10;
address_ina = 120;
address_inb = 121;
data_ina = 16'hb30;
data_inb = 16'h504;
#10;
address_ina = 122;
address_inb = 123;
data_ina = 16'h636;
data_inb = 16'h75a;
#10;
address_ina = 124;
address_inb = 125;
data_ina = 16'h7d9;
data_inb = 16'h18d;
#10;
address_ina = 126;
address_inb = 127;
data_ina = 16'h5d7;
data_inb = 16'h670;
#10;
address_ina = 128;
address_inb = 129;
data_ina = 16'h1c7;
data_inb = 16'h3b9;
#10;
address_ina = 130;
address_inb = 131;
data_ina = 16'ha4d;
data_inb = 16'h82a;
#10;
address_ina = 132;
address_inb = 133;
data_ina = 16'h81d;
data_inb = 16'h1e8;
#10;
address_ina = 134;
address_inb = 135;
data_ina = 16'hb19;
data_inb = 16'h135;
#10;
address_ina = 136;
address_inb = 137;
data_ina = 16'h246;
data_inb = 16'h60f;
#10;
address_ina = 138;
address_inb = 139;
data_ina = 16'h757;
data_inb = 16'h465;
#10;
address_ina = 140;
address_inb = 141;
data_ina = 16'hb10;
data_inb = 16'hbe0;
#10;
address_ina = 142;
address_inb = 143;
data_ina = 16'ha0c;
data_inb = 16'h56f;
#10;
address_ina = 144;
address_inb = 145;
data_ina = 16'hc03;
data_inb = 16'h914;
#10;
address_ina = 146;
address_inb = 147;
data_ina = 16'h858;
data_inb = 16'h4c0;
#10;
address_ina = 148;
address_inb = 149;
data_ina = 16'hac5;
data_inb = 16'ha02;
#10;
address_ina = 150;
address_inb = 151;
data_ina = 16'h72;
data_inb = 16'h5c4;
#10;
address_ina = 152;
address_inb = 153;
data_ina = 16'h650;
data_inb = 16'h9a3;
#10;
address_ina = 154;
address_inb = 155;
data_ina = 16'h336;
data_inb = 16'h259;
#10;
address_ina = 156;
address_inb = 157;
data_ina = 16'h747;
data_inb = 16'h434;
#10;
address_ina = 158;
address_inb = 159;
data_ina = 16'h78b;
data_inb = 16'h313;
#10;
address_ina = 160;
address_inb = 161;
data_ina = 16'h1aa;
data_inb = 16'h2b1;
#10;
address_ina = 162;
address_inb = 163;
data_ina = 16'h8d3;
data_inb = 16'h1fe;
#10;
address_ina = 164;
address_inb = 165;
data_ina = 16'hb06;
data_inb = 16'hc10;
#10;
address_ina = 166;
address_inb = 167;
data_ina = 16'hc7c;
data_inb = 16'h8b3;
#10;
address_ina = 168;
address_inb = 169;
data_ina = 16'h868;
data_inb = 16'h6d8;
#10;
address_ina = 170;
address_inb = 171;
data_ina = 16'hc9f;
data_inb = 16'h57c;
#10;
address_ina = 172;
address_inb = 173;
data_ina = 16'hcda;
data_inb = 16'h128;
#10;
address_ina = 174;
address_inb = 175;
data_ina = 16'h421;
data_inb = 16'h7f6;
#10;
address_ina = 176;
address_inb = 177;
data_ina = 16'he4;
data_inb = 16'h72d;
#10;
address_ina = 178;
address_inb = 179;
data_ina = 16'h8d7;
data_inb = 16'hd7;
#10;
address_ina = 180;
address_inb = 181;
data_ina = 16'h9e5;
data_inb = 16'h580;
#10;
address_ina = 182;
address_inb = 183;
data_ina = 16'hc96;
data_inb = 16'hc37;
#10;
address_ina = 184;
address_inb = 185;
data_ina = 16'hcf1;
data_inb = 16'h7ac;
#10;
address_ina = 186;
address_inb = 187;
data_ina = 16'h243;
data_inb = 16'h666;
#10;
address_ina = 188;
address_inb = 189;
data_ina = 16'h945;
data_inb = 16'h93f;
#10;
address_ina = 190;
address_inb = 191;
data_ina = 16'h862;
data_inb = 16'h1e1;
#10;
address_ina = 192;
address_inb = 193;
data_ina = 16'h22f;
data_inb = 16'h8d7;
#10;
address_ina = 194;
address_inb = 195;
data_ina = 16'hd;
data_inb = 16'hbd6;
#10;
address_ina = 196;
address_inb = 197;
data_ina = 16'hc2e;
data_inb = 16'hbbc;
#10;
address_ina = 198;
address_inb = 199;
data_ina = 16'hb57;
data_inb = 16'h11b;
#10;
address_ina = 200;
address_inb = 201;
data_ina = 16'hb5e;
data_inb = 16'h687;
#10;
address_ina = 202;
address_inb = 203;
data_ina = 16'h47f;
data_inb = 16'h771;
#10;
address_ina = 204;
address_inb = 205;
data_ina = 16'h8b9;
data_inb = 16'h892;
#10;
address_ina = 206;
address_inb = 207;
data_ina = 16'h225;
data_inb = 16'h18d;
#10;
address_ina = 208;
address_inb = 209;
data_ina = 16'h5fe;
data_inb = 16'h297;
#10;
address_ina = 210;
address_inb = 211;
data_ina = 16'h499;
data_inb = 16'hf1;
#10;
address_ina = 212;
address_inb = 213;
data_ina = 16'h186;
data_inb = 16'h2bb;
#10;
address_ina = 214;
address_inb = 215;
data_ina = 16'h656;
data_inb = 16'h559;
#10;
address_ina = 216;
address_inb = 217;
data_ina = 16'h4c0;
data_inb = 16'h3c2;
#10;
address_ina = 218;
address_inb = 219;
data_ina = 16'haf2;
data_inb = 16'h1e8;
#10;
address_ina = 220;
address_inb = 221;
data_ina = 16'h5d1;
data_inb = 16'h63f;
#10;
address_ina = 222;
address_inb = 223;
data_ina = 16'h889;
data_inb = 16'hadc;
#10;
address_ina = 224;
address_inb = 225;
data_ina = 16'h86b;
data_inb = 16'h51e;
#10;
address_ina = 226;
address_inb = 227;
data_ina = 16'ha33;
data_inb = 16'h8c;
#10;
address_ina = 228;
address_inb = 229;
data_ina = 16'h4f4;
data_inb = 16'h46f;
#10;
address_ina = 230;
address_inb = 231;
data_ina = 16'hb40;
data_inb = 16'ha91;
#10;
address_ina = 232;
address_inb = 233;
data_ina = 16'h94f;
data_inb = 16'h4c6;
#10;
address_ina = 234;
address_inb = 235;
data_ina = 16'h212;
data_inb = 16'ha9b;
#10;
address_ina = 236;
address_inb = 237;
data_ina = 16'had5;
data_inb = 16'ha3c;
#10;
address_ina = 238;
address_inb = 239;
data_ina = 16'h14c;
data_inb = 16'h639;
#10;
address_ina = 240;
address_inb = 241;
data_ina = 16'h21c;
data_inb = 16'h28d;
#10;
address_ina = 242;
address_inb = 243;
data_ina = 16'h576;
data_inb = 16'hb85;
#10;
address_ina = 244;
address_inb = 245;
data_ina = 16'hacb;
data_inb = 16'h966;
#10;
address_ina = 246;
address_inb = 247;
data_ina = 16'h8d3;
data_inb = 16'h555;
#10;
address_ina = 248;
address_inb = 249;
data_ina = 16'h3fd;
data_inb = 16'ha2c;
#10;
address_ina = 250;
address_inb = 251;
data_ina = 16'h82;
data_inb = 16'h681;
#10;
address_ina = 252;
address_inb = 253;
data_ina = 16'haec;
data_inb = 16'h744;
#10;
address_ina = 254;
address_inb = 255;
data_ina = 16'hcd7;
data_inb = 16'h259;
#10;
        wait(init_done);
        #30
        we = 0;
        // Start processing
         
		  #38000

        start = 0;



//        wait (wr_req);
//		  wait (!wr_req);
//		   rd_req = 1;
		  wait(done);
		  #20000
rd_req = 1;
        #70 
		  start = 1;
		 #80 
wait(rd_empty)
rd_req = 0;

$display("Finished the NTT test Number %d",test_num);
////Begin test number #44//////////////
rst = 1;

//#1000
start = 1;
mode = 0; //NTT 0 // INTT 1

// Reset for a few clock cycles

#1000

rst = 0;
test_num = test_num + 1;
#1000
we = 1;
address_ina = 0;
address_inb = 1;
data_ina = 16'h344;
data_inb = 16'hcf7;
#10;
address_ina = 2;
address_inb = 3;
data_ina = 16'h37e;
data_inb = 16'ha70;
#10;
address_ina = 4;
address_inb = 5;
data_ina = 16'h996;
data_inb = 16'h862;
#10;
address_ina = 6;
address_inb = 7;
data_ina = 16'ha5d;
data_inb = 16'h20f;
#10;
address_ina = 8;
address_inb = 9;
data_ina = 16'h125;
data_inb = 16'h8a3;
#10;
address_ina = 10;
address_inb = 11;
data_ina = 16'h824;
data_inb = 16'h17;
#10;
address_ina = 12;
address_inb = 13;
data_ina = 16'h3f3;
data_inb = 16'h615;
#10;
address_ina = 14;
address_inb = 15;
data_ina = 16'h263;
data_inb = 16'hcac;
#10;
address_ina = 16;
address_inb = 17;
data_ina = 16'h340;
data_inb = 16'h70c;
#10;
address_ina = 18;
address_inb = 19;
data_ina = 16'h59d;
data_inb = 16'h9ad;
#10;
address_ina = 20;
address_inb = 21;
data_ina = 16'h8f;
data_inb = 16'h8a6;
#10;
address_ina = 22;
address_inb = 23;
data_ina = 16'hb7e;
data_inb = 16'h593;
#10;
address_ina = 24;
address_inb = 25;
data_ina = 16'h1c7;
data_inb = 16'h865;
#10;
address_ina = 26;
address_inb = 27;
data_ina = 16'h388;
data_inb = 16'h482;
#10;
address_ina = 28;
address_inb = 29;
data_ina = 16'h629;
data_inb = 16'h61f;
#10;
address_ina = 30;
address_inb = 31;
data_ina = 16'h3e6;
data_inb = 16'h18d;
#10;
address_ina = 32;
address_inb = 33;
data_ina = 16'h841;
data_inb = 16'h1e4;
#10;
address_ina = 34;
address_inb = 35;
data_ina = 16'hbd;
data_inb = 16'h400;
#10;
address_ina = 36;
address_inb = 37;
data_ina = 16'ha1f;
data_inb = 16'h942;
#10;
address_ina = 38;
address_inb = 39;
data_ina = 16'h2b1;
data_inb = 16'h862;
#10;
address_ina = 40;
address_inb = 41;
data_ina = 16'h1e4;
data_inb = 16'hb6;
#10;
address_ina = 42;
address_inb = 43;
data_ina = 16'h36b;
data_inb = 16'h821;
#10;
address_ina = 44;
address_inb = 45;
data_ina = 16'hd3;
data_inb = 16'ha6;
#10;
address_ina = 46;
address_inb = 47;
data_ina = 16'hc5e;
data_inb = 16'hc96;
#10;
address_ina = 48;
address_inb = 49;
data_ina = 16'h46b;
data_inb = 16'ha5d;
#10;
address_ina = 50;
address_inb = 51;
data_ina = 16'hc0;
data_inb = 16'h504;
#10;
address_ina = 52;
address_inb = 53;
data_ina = 16'h656;
data_inb = 16'h441;
#10;
address_ina = 54;
address_inb = 55;
data_ina = 16'ha4d;
data_inb = 16'h53b;
#10;
address_ina = 56;
address_inb = 57;
data_ina = 16'h65d;
data_inb = 16'h1b7;
#10;
address_ina = 58;
address_inb = 59;
data_ina = 16'h62;
data_inb = 16'h583;
#10;
address_ina = 60;
address_inb = 61;
data_ina = 16'hb2a;
data_inb = 16'h3f3;
#10;
address_ina = 62;
address_inb = 63;
data_ina = 16'h492;
data_inb = 16'h196;
#10;
address_ina = 64;
address_inb = 65;
data_ina = 16'h326;
data_inb = 16'ha70;
#10;
address_ina = 66;
address_inb = 67;
data_ina = 16'hcfa;
data_inb = 16'h7bc;
#10;
address_ina = 68;
address_inb = 69;
data_ina = 16'h15f;
data_inb = 16'h938;
#10;
address_ina = 70;
address_inb = 71;
data_ina = 16'h492;
data_inb = 16'hb3a;
#10;
address_ina = 72;
address_inb = 73;
data_ina = 16'h5eb;
data_inb = 16'h395;
#10;
address_ina = 74;
address_inb = 75;
data_ina = 16'hc37;
data_inb = 16'hb57;
#10;
address_ina = 76;
address_inb = 77;
data_ina = 16'hb7b;
data_inb = 16'h72d;
#10;
address_ina = 78;
address_inb = 79;
data_ina = 16'h62f;
data_inb = 16'h71d;
#10;
address_ina = 80;
address_inb = 81;
data_ina = 16'h33d;
data_inb = 16'h89f;
#10;
address_ina = 82;
address_inb = 83;
data_ina = 16'h50e;
data_inb = 16'h1ce;
#10;
address_ina = 84;
address_inb = 85;
data_ina = 16'h6f9;
data_inb = 16'h9c;
#10;
address_ina = 86;
address_inb = 87;
data_ina = 16'h792;
data_inb = 16'h378;
#10;
address_ina = 88;
address_inb = 89;
data_ina = 16'h431;
data_inb = 16'ha29;
#10;
address_ina = 90;
address_inb = 91;
data_ina = 16'h3e6;
data_inb = 16'h8e0;
#10;
address_ina = 92;
address_inb = 93;
data_ina = 16'h691;
data_inb = 16'hc6f;
#10;
address_ina = 94;
address_inb = 95;
data_ina = 16'hb9;
data_inb = 16'h6d5;
#10;
address_ina = 96;
address_inb = 97;
data_ina = 16'h7b9;
data_inb = 16'h51;
#10;
address_ina = 98;
address_inb = 99;
data_ina = 16'ha91;
data_inb = 16'h548;
#10;
address_ina = 100;
address_inb = 101;
data_ina = 16'ha1c;
data_inb = 16'h2ec;
#10;
address_ina = 102;
address_inb = 103;
data_ina = 16'h11e;
data_inb = 16'hc8c;
#10;
address_ina = 104;
address_inb = 105;
data_ina = 16'h7b9;
data_inb = 16'h132;
#10;
address_ina = 106;
address_inb = 107;
data_ina = 16'h2b8;
data_inb = 16'h9ff;
#10;
address_ina = 108;
address_inb = 109;
data_ina = 16'h91b;
data_inb = 16'h82a;
#10;
address_ina = 110;
address_inb = 111;
data_ina = 16'h844;
data_inb = 16'h499;
#10;
address_ina = 112;
address_inb = 113;
data_ina = 16'hcbd;
data_inb = 16'h427;
#10;
address_ina = 114;
address_inb = 115;
data_ina = 16'h61f;
data_inb = 16'h8c;
#10;
address_ina = 116;
address_inb = 117;
data_ina = 16'hcfe;
data_inb = 16'h2db;
#10;
address_ina = 118;
address_inb = 119;
data_ina = 16'ha84;
data_inb = 16'h4f4;
#10;
address_ina = 120;
address_inb = 121;
data_ina = 16'h492;
data_inb = 16'h899;
#10;
address_ina = 122;
address_inb = 123;
data_ina = 16'h9ce;
data_inb = 16'h2d2;
#10;
address_ina = 124;
address_inb = 125;
data_ina = 16'h962;
data_inb = 16'h86b;
#10;
address_ina = 126;
address_inb = 127;
data_ina = 16'h42a;
data_inb = 16'h25d;
#10;
address_ina = 128;
address_inb = 129;
data_ina = 16'h54f;
data_inb = 16'hb64;
#10;
address_ina = 130;
address_inb = 131;
data_ina = 16'h781;
data_inb = 16'h9cb;
#10;
address_ina = 132;
address_inb = 133;
data_ina = 16'h1fb;
data_inb = 16'h5b0;
#10;
address_ina = 134;
address_inb = 135;
data_ina = 16'h54c;
data_inb = 16'h6ae;
#10;
address_ina = 136;
address_inb = 137;
data_ina = 16'h7b9;
data_inb = 16'h186;
#10;
address_ina = 138;
address_inb = 139;
data_ina = 16'h388;
data_inb = 16'h3c6;
#10;
address_ina = 140;
address_inb = 141;
data_ina = 16'h14c;
data_inb = 16'h5b0;
#10;
address_ina = 142;
address_inb = 143;
data_ina = 16'hc51;
data_inb = 16'ha9e;
#10;
address_ina = 144;
address_inb = 145;
data_ina = 16'h9a7;
data_inb = 16'hb44;
#10;
address_ina = 146;
address_inb = 147;
data_ina = 16'h96f;
data_inb = 16'ha7a;
#10;
address_ina = 148;
address_inb = 149;
data_ina = 16'h478;
data_inb = 16'h496;
#10;
address_ina = 150;
address_inb = 151;
data_ina = 16'h7d3;
data_inb = 16'h92e;
#10;
address_ina = 152;
address_inb = 153;
data_ina = 16'h61f;
data_inb = 16'h2ab;
#10;
address_ina = 154;
address_inb = 155;
data_ina = 16'h73a;
data_inb = 16'hbe6;
#10;
address_ina = 156;
address_inb = 157;
data_ina = 16'hbfd;
data_inb = 16'h421;
#10;
address_ina = 158;
address_inb = 159;
data_ina = 16'h44b;
data_inb = 16'h8b6;
#10;
address_ina = 160;
address_inb = 161;
data_ina = 16'h7bc;
data_inb = 16'h5c4;
#10;
address_ina = 162;
address_inb = 163;
data_ina = 16'h8b6;
data_inb = 16'h774;
#10;
address_ina = 164;
address_inb = 165;
data_ina = 16'h4a9;
data_inb = 16'h169;
#10;
address_ina = 166;
address_inb = 167;
data_ina = 16'h885;
data_inb = 16'hb16;
#10;
address_ina = 168;
address_inb = 169;
data_ina = 16'h259;
data_inb = 16'h740;
#10;
address_ina = 170;
address_inb = 171;
data_ina = 16'h778;
data_inb = 16'hab1;
#10;
address_ina = 172;
address_inb = 173;
data_ina = 16'h875;
data_inb = 16'hd0;
#10;
address_ina = 174;
address_inb = 175;
data_ina = 16'hb0;
data_inb = 16'h4b;
#10;
address_ina = 176;
address_inb = 177;
data_ina = 16'h865;
data_inb = 16'h980;
#10;
address_ina = 178;
address_inb = 179;
data_ina = 16'h3d3;
data_inb = 16'habb;
#10;
address_ina = 180;
address_inb = 181;
data_ina = 16'h410;
data_inb = 16'ha3c;
#10;
address_ina = 182;
address_inb = 183;
data_ina = 16'h69b;
data_inb = 16'hac5;
#10;
address_ina = 184;
address_inb = 185;
data_ina = 16'h97c;
data_inb = 16'h834;
#10;
address_ina = 186;
address_inb = 187;
data_ina = 16'ha8a;
data_inb = 16'h266;
#10;
address_ina = 188;
address_inb = 189;
data_ina = 16'hb7b;
data_inb = 16'h5f8;
#10;
address_ina = 190;
address_inb = 191;
data_ina = 16'h4ca;
data_inb = 16'hac2;
#10;
address_ina = 192;
address_inb = 193;
data_ina = 16'h72a;
data_inb = 16'h878;
#10;
address_ina = 194;
address_inb = 195;
data_ina = 16'h1e1;
data_inb = 16'h7af;
#10;
address_ina = 196;
address_inb = 197;
data_ina = 16'h11b;
data_inb = 16'h596;
#10;
address_ina = 198;
address_inb = 199;
data_ina = 16'hca;
data_inb = 16'h6a4;
#10;
address_ina = 200;
address_inb = 201;
data_ina = 16'hb09;
data_inb = 16'h996;
#10;
address_ina = 202;
address_inb = 203;
data_ina = 16'h8fa;
data_inb = 16'h7fa;
#10;
address_ina = 204;
address_inb = 205;
data_ina = 16'h83b;
data_inb = 16'h730;
#10;
address_ina = 206;
address_inb = 207;
data_ina = 16'h3e0;
data_inb = 16'h448;
#10;
address_ina = 208;
address_inb = 209;
data_ina = 16'h7f3;
data_inb = 16'h1c7;
#10;
address_ina = 210;
address_inb = 211;
data_ina = 16'h911;
data_inb = 16'hc5b;
#10;
address_ina = 212;
address_inb = 213;
data_ina = 16'h990;
data_inb = 16'h1c7;
#10;
address_ina = 214;
address_inb = 215;
data_ina = 16'hb1d;
data_inb = 16'ha0c;
#10;
address_ina = 216;
address_inb = 217;
data_ina = 16'ha4d;
data_inb = 16'h538;
#10;
address_ina = 218;
address_inb = 219;
data_ina = 16'hbe9;
data_inb = 16'h9bd;
#10;
address_ina = 220;
address_inb = 221;
data_ina = 16'h636;
data_inb = 16'hbe6;
#10;
address_ina = 222;
address_inb = 223;
data_ina = 16'h2b4;
data_inb = 16'h38e;
#10;
address_ina = 224;
address_inb = 225;
data_ina = 16'hbdc;
data_inb = 16'hb3d;
#10;
address_ina = 226;
address_inb = 227;
data_ina = 16'h319;
data_inb = 16'hca6;
#10;
address_ina = 228;
address_inb = 229;
data_ina = 16'h118;
data_inb = 16'h8d0;
#10;
address_ina = 230;
address_inb = 231;
data_ina = 16'h6be;
data_inb = 16'h56f;
#10;
address_ina = 232;
address_inb = 233;
data_ina = 16'h4a3;
data_inb = 16'h7bc;
#10;
address_ina = 234;
address_inb = 235;
data_ina = 16'h51e;
data_inb = 16'h27;
#10;
address_ina = 236;
address_inb = 237;
data_ina = 16'h8da;
data_inb = 16'h4a9;
#10;
address_ina = 238;
address_inb = 239;
data_ina = 16'h9cb;
data_inb = 16'h13b;
#10;
address_ina = 240;
address_inb = 241;
data_ina = 16'h608;
data_inb = 16'h55f;
#10;
address_ina = 242;
address_inb = 243;
data_ina = 16'h3d3;
data_inb = 16'hb51;
#10;
address_ina = 244;
address_inb = 245;
data_ina = 16'hb10;
data_inb = 16'h5f5;
#10;
address_ina = 246;
address_inb = 247;
data_ina = 16'h57c;
data_inb = 16'h4e;
#10;
address_ina = 248;
address_inb = 249;
data_ina = 16'h744;
data_inb = 16'h573;
#10;
address_ina = 250;
address_inb = 251;
data_ina = 16'h4c6;
data_inb = 16'hc7f;
#10;
address_ina = 252;
address_inb = 253;
data_ina = 16'h5c7;
data_inb = 16'h51e;
#10;
address_ina = 254;
address_inb = 255;
data_ina = 16'hcd3;
data_inb = 16'h193;
#10;
        wait(init_done);
        #30
        we = 0;
        // Start processing
         
		  #38000

        start = 0;



//        wait (wr_req);
//		  wait (!wr_req);
//		   rd_req = 1;
		  wait(done);
		  #20000
rd_req = 1;
        #70 
		  start = 1;
		 #80 
wait(rd_empty)
rd_req = 0;

$display("Finished the NTT test Number %d",test_num);
////Begin test number #45//////////////
rst = 1;

//#1000
start = 1;
mode = 1; //NTT 0 // INTT 1

// Reset for a few clock cycles

#1000

rst = 0;
test_num = test_num + 1;
#1000
we = 1;
address_ina = 0;
address_inb = 1;
data_ina = 16'h2b4;
data_inb = 16'hf9fb;
#10;
address_ina = 2;
address_inb = 3;
data_ina = 16'h41d;
data_inb = 16'hfa06;
#10;
address_ina = 4;
address_inb = 5;
data_ina = 16'hfebc;
data_inb = 16'hfc49;
#10;
address_ina = 6;
address_inb = 7;
data_ina = 16'hfb27;
data_inb = 16'hfde2;
#10;
address_ina = 8;
address_inb = 9;
data_ina = 16'h5a3;
data_inb = 16'hfde7;
#10;
address_ina = 10;
address_inb = 11;
data_ina = 16'h1d0;
data_inb = 16'hfa92;
#10;
address_ina = 12;
address_inb = 13;
data_ina = 16'h1c1;
data_inb = 16'hfd66;
#10;
address_ina = 14;
address_inb = 15;
data_ina = 16'h124;
data_inb = 16'hfd8a;
#10;
address_ina = 16;
address_inb = 17;
data_ina = 16'hfc80;
data_inb = 16'h392;
#10;
address_ina = 18;
address_inb = 19;
data_ina = 16'hffd8;
data_inb = 16'hfa16;
#10;
address_ina = 20;
address_inb = 21;
data_ina = 16'hfbf7;
data_inb = 16'hfed5;
#10;
address_ina = 22;
address_inb = 23;
data_ina = 16'hfc7e;
data_inb = 16'hf9eb;
#10;
address_ina = 24;
address_inb = 25;
data_ina = 16'h113;
data_inb = 16'hf989;
#10;
address_ina = 26;
address_inb = 27;
data_ina = 16'h264;
data_inb = 16'hfae7;
#10;
address_ina = 28;
address_inb = 29;
data_ina = 16'hfc54;
data_inb = 16'h565;
#10;
address_ina = 30;
address_inb = 31;
data_ina = 16'hfa6a;
data_inb = 16'h10c;
#10;
address_ina = 32;
address_inb = 33;
data_ina = 16'h4ae;
data_inb = 16'h3e;
#10;
address_ina = 34;
address_inb = 35;
data_ina = 16'h3f9;
data_inb = 16'hfb10;
#10;
address_ina = 36;
address_inb = 37;
data_ina = 16'h372;
data_inb = 16'hfaa3;
#10;
address_ina = 38;
address_inb = 39;
data_ina = 16'h511;
data_inb = 16'hfc26;
#10;
address_ina = 40;
address_inb = 41;
data_ina = 16'hfe08;
data_inb = 16'hfff2;
#10;
address_ina = 42;
address_inb = 43;
data_ina = 16'h1a3;
data_inb = 16'h20b;
#10;
address_ina = 44;
address_inb = 45;
data_ina = 16'hc9;
data_inb = 16'hc0;
#10;
address_ina = 46;
address_inb = 47;
data_ina = 16'h5b4;
data_inb = 16'hfa1b;
#10;
address_ina = 48;
address_inb = 49;
data_ina = 16'h640;
data_inb = 16'h4a;
#10;
address_ina = 50;
address_inb = 51;
data_ina = 16'h423;
data_inb = 16'h4f2;
#10;
address_ina = 52;
address_inb = 53;
data_ina = 16'hfa55;
data_inb = 16'h2bd;
#10;
address_ina = 54;
address_inb = 55;
data_ina = 16'h150;
data_inb = 16'h31a;
#10;
address_ina = 56;
address_inb = 57;
data_ina = 16'h31b;
data_inb = 16'hfcd7;
#10;
address_ina = 58;
address_inb = 59;
data_ina = 16'h278;
data_inb = 16'h54e;
#10;
address_ina = 60;
address_inb = 61;
data_ina = 16'hfc5b;
data_inb = 16'hfff3;
#10;
address_ina = 62;
address_inb = 63;
data_ina = 16'h5ee;
data_inb = 16'hfdaf;
#10;
address_ina = 64;
address_inb = 65;
data_ina = 16'hffbe;
data_inb = 16'hf9be;
#10;
address_ina = 66;
address_inb = 67;
data_ina = 16'h49d;
data_inb = 16'h34b;
#10;
address_ina = 68;
address_inb = 69;
data_ina = 16'h102;
data_inb = 16'h50a;
#10;
address_ina = 70;
address_inb = 71;
data_ina = 16'hfb64;
data_inb = 16'h0;
#10;
address_ina = 72;
address_inb = 73;
data_ina = 16'h219;
data_inb = 16'h224;
#10;
address_ina = 74;
address_inb = 75;
data_ina = 16'h41;
data_inb = 16'h2e9;
#10;
address_ina = 76;
address_inb = 77;
data_ina = 16'hfc6a;
data_inb = 16'hfa7c;
#10;
address_ina = 78;
address_inb = 79;
data_ina = 16'hfd4f;
data_inb = 16'h54c;
#10;
address_ina = 80;
address_inb = 81;
data_ina = 16'h97;
data_inb = 16'hfca4;
#10;
address_ina = 82;
address_inb = 83;
data_ina = 16'hfcac;
data_inb = 16'hfa69;
#10;
address_ina = 84;
address_inb = 85;
data_ina = 16'hf9c0;
data_inb = 16'h29e;
#10;
address_ina = 86;
address_inb = 87;
data_ina = 16'hff87;
data_inb = 16'hf9cb;
#10;
address_ina = 88;
address_inb = 89;
data_ina = 16'h25c;
data_inb = 16'h4da;
#10;
address_ina = 90;
address_inb = 91;
data_ina = 16'hfb37;
data_inb = 16'h26e;
#10;
address_ina = 92;
address_inb = 93;
data_ina = 16'hfc5d;
data_inb = 16'hfad8;
#10;
address_ina = 94;
address_inb = 95;
data_ina = 16'hffef;
data_inb = 16'hfb4e;
#10;
address_ina = 96;
address_inb = 97;
data_ina = 16'hfa7c;
data_inb = 16'h633;
#10;
address_ina = 98;
address_inb = 99;
data_ina = 16'hdb;
data_inb = 16'hfdaf;
#10;
address_ina = 100;
address_inb = 101;
data_ina = 16'h530;
data_inb = 16'hf9c7;
#10;
address_ina = 102;
address_inb = 103;
data_ina = 16'hf9f6;
data_inb = 16'h29f;
#10;
address_ina = 104;
address_inb = 105;
data_ina = 16'hf994;
data_inb = 16'hf9ea;
#10;
address_ina = 106;
address_inb = 107;
data_ina = 16'hfc59;
data_inb = 16'hfefd;
#10;
address_ina = 108;
address_inb = 109;
data_ina = 16'hfd85;
data_inb = 16'h4c0;
#10;
address_ina = 110;
address_inb = 111;
data_ina = 16'hfd58;
data_inb = 16'hfeda;
#10;
address_ina = 112;
address_inb = 113;
data_ina = 16'hf9af;
data_inb = 16'hfa58;
#10;
address_ina = 114;
address_inb = 115;
data_ina = 16'h30a;
data_inb = 16'h65e;
#10;
address_ina = 116;
address_inb = 117;
data_ina = 16'h303;
data_inb = 16'hf9c7;
#10;
address_ina = 118;
address_inb = 119;
data_ina = 16'hfb2d;
data_inb = 16'h503;
#10;
address_ina = 120;
address_inb = 121;
data_ina = 16'hfdd0;
data_inb = 16'hfee4;
#10;
address_ina = 122;
address_inb = 123;
data_ina = 16'h202;
data_inb = 16'hff59;
#10;
address_ina = 124;
address_inb = 125;
data_ina = 16'h2c9;
data_inb = 16'h30b;
#10;
address_ina = 126;
address_inb = 127;
data_ina = 16'h4e3;
data_inb = 16'hff9b;
#10;
address_ina = 128;
address_inb = 129;
data_ina = 16'hfcad;
data_inb = 16'hfa6f;
#10;
address_ina = 130;
address_inb = 131;
data_ina = 16'hffc6;
data_inb = 16'hfdad;
#10;
address_ina = 132;
address_inb = 133;
data_ina = 16'h40e;
data_inb = 16'h4fd;
#10;
address_ina = 134;
address_inb = 135;
data_ina = 16'hfef1;
data_inb = 16'h66e;
#10;
address_ina = 136;
address_inb = 137;
data_ina = 16'h28c;
data_inb = 16'hfac8;
#10;
address_ina = 138;
address_inb = 139;
data_ina = 16'hffdd;
data_inb = 16'hf9a9;
#10;
address_ina = 140;
address_inb = 141;
data_ina = 16'hfa98;
data_inb = 16'h28d;
#10;
address_ina = 142;
address_inb = 143;
data_ina = 16'h35b;
data_inb = 16'hfb98;
#10;
address_ina = 144;
address_inb = 145;
data_ina = 16'h486;
data_inb = 16'hffa5;
#10;
address_ina = 146;
address_inb = 147;
data_ina = 16'hfcde;
data_inb = 16'h4ae;
#10;
address_ina = 148;
address_inb = 149;
data_ina = 16'h244;
data_inb = 16'hfb7f;
#10;
address_ina = 150;
address_inb = 151;
data_ina = 16'h4be;
data_inb = 16'h2f2;
#10;
address_ina = 152;
address_inb = 153;
data_ina = 16'h127;
data_inb = 16'hfe49;
#10;
address_ina = 154;
address_inb = 155;
data_ina = 16'h2df;
data_inb = 16'h57f;
#10;
address_ina = 156;
address_inb = 157;
data_ina = 16'h264;
data_inb = 16'hdd;
#10;
address_ina = 158;
address_inb = 159;
data_ina = 16'hfc3d;
data_inb = 16'h579;
#10;
address_ina = 160;
address_inb = 161;
data_ina = 16'h4bc;
data_inb = 16'hfacb;
#10;
address_ina = 162;
address_inb = 163;
data_ina = 16'hfb36;
data_inb = 16'hfbba;
#10;
address_ina = 164;
address_inb = 165;
data_ina = 16'hff88;
data_inb = 16'h3f3;
#10;
address_ina = 166;
address_inb = 167;
data_ina = 16'h38b;
data_inb = 16'h2ac;
#10;
address_ina = 168;
address_inb = 169;
data_ina = 16'hfa2d;
data_inb = 16'hf0;
#10;
address_ina = 170;
address_inb = 171;
data_ina = 16'h3aa;
data_inb = 16'h113;
#10;
address_ina = 172;
address_inb = 173;
data_ina = 16'hfcca;
data_inb = 16'hfcc3;
#10;
address_ina = 174;
address_inb = 175;
data_ina = 16'h47a;
data_inb = 16'h4d5;
#10;
address_ina = 176;
address_inb = 177;
data_ina = 16'h2ba;
data_inb = 16'h405;
#10;
address_ina = 178;
address_inb = 179;
data_ina = 16'h3b1;
data_inb = 16'hfc14;
#10;
address_ina = 180;
address_inb = 181;
data_ina = 16'hfd8b;
data_inb = 16'hfdaa;
#10;
address_ina = 182;
address_inb = 183;
data_ina = 16'hfae7;
data_inb = 16'hb5;
#10;
address_ina = 184;
address_inb = 185;
data_ina = 16'hffa0;
data_inb = 16'hfa7d;
#10;
address_ina = 186;
address_inb = 187;
data_ina = 16'h1e8;
data_inb = 16'hb7;
#10;
address_ina = 188;
address_inb = 189;
data_ina = 16'h242;
data_inb = 16'hf9a2;
#10;
address_ina = 190;
address_inb = 191;
data_ina = 16'hfe9e;
data_inb = 16'h3b4;
#10;
address_ina = 192;
address_inb = 193;
data_ina = 16'h453;
data_inb = 16'h127;
#10;
address_ina = 194;
address_inb = 195;
data_ina = 16'h2b7;
data_inb = 16'h62e;
#10;
address_ina = 196;
address_inb = 197;
data_ina = 16'h1a0;
data_inb = 16'h55c;
#10;
address_ina = 198;
address_inb = 199;
data_ina = 16'hfd8a;
data_inb = 16'h161;
#10;
address_ina = 200;
address_inb = 201;
data_ina = 16'hfd34;
data_inb = 16'hfc9e;
#10;
address_ina = 202;
address_inb = 203;
data_ina = 16'hfa27;
data_inb = 16'hfc97;
#10;
address_ina = 204;
address_inb = 205;
data_ina = 16'h3c9;
data_inb = 16'hfe5f;
#10;
address_ina = 206;
address_inb = 207;
data_ina = 16'hfde6;
data_inb = 16'hffd3;
#10;
address_ina = 208;
address_inb = 209;
data_ina = 16'h223;
data_inb = 16'hfd98;
#10;
address_ina = 210;
address_inb = 211;
data_ina = 16'hff7e;
data_inb = 16'hfa2a;
#10;
address_ina = 212;
address_inb = 213;
data_ina = 16'hffd2;
data_inb = 16'h602;
#10;
address_ina = 214;
address_inb = 215;
data_ina = 16'h15d;
data_inb = 16'hfbef;
#10;
address_ina = 216;
address_inb = 217;
data_ina = 16'hfb11;
data_inb = 16'h55e;
#10;
address_ina = 218;
address_inb = 219;
data_ina = 16'h1bb;
data_inb = 16'h10d;
#10;
address_ina = 220;
address_inb = 221;
data_ina = 16'hfdb6;
data_inb = 16'hfb11;
#10;
address_ina = 222;
address_inb = 223;
data_ina = 16'h49b;
data_inb = 16'hfc0e;
#10;
address_ina = 224;
address_inb = 225;
data_ina = 16'h41;
data_inb = 16'h26;
#10;
address_ina = 226;
address_inb = 227;
data_ina = 16'h196;
data_inb = 16'hfa63;
#10;
address_ina = 228;
address_inb = 229;
data_ina = 16'h2b;
data_inb = 16'hfaf6;
#10;
address_ina = 230;
address_inb = 231;
data_ina = 16'hfd45;
data_inb = 16'hfb9a;
#10;
address_ina = 232;
address_inb = 233;
data_ina = 16'h2b6;
data_inb = 16'hfc74;
#10;
address_ina = 234;
address_inb = 235;
data_ina = 16'h5c9;
data_inb = 16'hfc27;
#10;
address_ina = 236;
address_inb = 237;
data_ina = 16'hf9af;
data_inb = 16'h148;
#10;
address_ina = 238;
address_inb = 239;
data_ina = 16'h358;
data_inb = 16'hfbf9;
#10;
address_ina = 240;
address_inb = 241;
data_ina = 16'h49a;
data_inb = 16'hfa93;
#10;
address_ina = 242;
address_inb = 243;
data_ina = 16'hfeba;
data_inb = 16'hfa02;
#10;
address_ina = 244;
address_inb = 245;
data_ina = 16'hfca2;
data_inb = 16'heb;
#10;
address_ina = 246;
address_inb = 247;
data_ina = 16'hff30;
data_inb = 16'hfd23;
#10;
address_ina = 248;
address_inb = 249;
data_ina = 16'h649;
data_inb = 16'h412;
#10;
address_ina = 250;
address_inb = 251;
data_ina = 16'hff0a;
data_inb = 16'h3ab;
#10;
address_ina = 252;
address_inb = 253;
data_ina = 16'hfabb;
data_inb = 16'h49f;
#10;
address_ina = 254;
address_inb = 255;
data_ina = 16'hfd85;
data_inb = 16'hfe66;
#10;
        wait(init_done);
        #30
        we = 0;
        // Start processing
         
		  #38000

        start = 0;



//        wait (wr_req);
//		  wait (!wr_req);
//		   rd_req = 1;
		  wait(done);
		  #20000
rd_req = 1;
        #70 
		  start = 1;
		 #80 
wait(rd_empty)
rd_req = 0;

$display("Finished the NTT test Number %d",test_num);
////Begin test number #46//////////////
rst = 1;

//#1000
start = 1;
mode = 0; //NTT 0 // INTT 1

// Reset for a few clock cycles

#1000

rst = 0;
test_num = test_num + 1;
#1000
we = 1;
address_ina = 0;
address_inb = 1;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 2;
address_inb = 3;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 4;
address_inb = 5;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 6;
address_inb = 7;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 8;
address_inb = 9;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 10;
address_inb = 11;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 12;
address_inb = 13;
data_ina = 16'h0;
data_inb = 16'h2;
#10;
address_ina = 14;
address_inb = 15;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 16;
address_inb = 17;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 18;
address_inb = 19;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 20;
address_inb = 21;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 22;
address_inb = 23;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 24;
address_inb = 25;
data_ina = 16'hfffe;
data_inb = 16'hfffe;
#10;
address_ina = 26;
address_inb = 27;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 28;
address_inb = 29;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 30;
address_inb = 31;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 32;
address_inb = 33;
data_ina = 16'h0;
data_inb = 16'h2;
#10;
address_ina = 34;
address_inb = 35;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 36;
address_inb = 37;
data_ina = 16'h1;
data_inb = 16'hfffe;
#10;
address_ina = 38;
address_inb = 39;
data_ina = 16'h2;
data_inb = 16'hfffe;
#10;
address_ina = 40;
address_inb = 41;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 42;
address_inb = 43;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 44;
address_inb = 45;
data_ina = 16'h0;
data_inb = 16'h2;
#10;
address_ina = 46;
address_inb = 47;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 48;
address_inb = 49;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 50;
address_inb = 51;
data_ina = 16'hfffe;
data_inb = 16'h0;
#10;
address_ina = 52;
address_inb = 53;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 54;
address_inb = 55;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 56;
address_inb = 57;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 58;
address_inb = 59;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 60;
address_inb = 61;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 62;
address_inb = 63;
data_ina = 16'h2;
data_inb = 16'hffff;
#10;
address_ina = 64;
address_inb = 65;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 66;
address_inb = 67;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 68;
address_inb = 69;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 70;
address_inb = 71;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 72;
address_inb = 73;
data_ina = 16'hffff;
data_inb = 16'hfffe;
#10;
address_ina = 74;
address_inb = 75;
data_ina = 16'h2;
data_inb = 16'h0;
#10;
address_ina = 76;
address_inb = 77;
data_ina = 16'hffff;
data_inb = 16'h2;
#10;
address_ina = 78;
address_inb = 79;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 80;
address_inb = 81;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 82;
address_inb = 83;
data_ina = 16'h2;
data_inb = 16'h0;
#10;
address_ina = 84;
address_inb = 85;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 86;
address_inb = 87;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 88;
address_inb = 89;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 90;
address_inb = 91;
data_ina = 16'hffff;
data_inb = 16'hfffe;
#10;
address_ina = 92;
address_inb = 93;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 94;
address_inb = 95;
data_ina = 16'h2;
data_inb = 16'h1;
#10;
address_ina = 96;
address_inb = 97;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 98;
address_inb = 99;
data_ina = 16'h0;
data_inb = 16'h2;
#10;
address_ina = 100;
address_inb = 101;
data_ina = 16'h0;
data_inb = 16'hfffe;
#10;
address_ina = 102;
address_inb = 103;
data_ina = 16'h2;
data_inb = 16'h0;
#10;
address_ina = 104;
address_inb = 105;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 106;
address_inb = 107;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 108;
address_inb = 109;
data_ina = 16'hfffe;
data_inb = 16'hffff;
#10;
address_ina = 110;
address_inb = 111;
data_ina = 16'hfffd;
data_inb = 16'h1;
#10;
address_ina = 112;
address_inb = 113;
data_ina = 16'h0;
data_inb = 16'hfffe;
#10;
address_ina = 114;
address_inb = 115;
data_ina = 16'hfffe;
data_inb = 16'hfffe;
#10;
address_ina = 116;
address_inb = 117;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 118;
address_inb = 119;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 120;
address_inb = 121;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 122;
address_inb = 123;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 124;
address_inb = 125;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 126;
address_inb = 127;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 128;
address_inb = 129;
data_ina = 16'h2;
data_inb = 16'hfffd;
#10;
address_ina = 130;
address_inb = 131;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 132;
address_inb = 133;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 134;
address_inb = 135;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 136;
address_inb = 137;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 138;
address_inb = 139;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 140;
address_inb = 141;
data_ina = 16'h0;
data_inb = 16'h2;
#10;
address_ina = 142;
address_inb = 143;
data_ina = 16'hfffd;
data_inb = 16'h0;
#10;
address_ina = 144;
address_inb = 145;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 146;
address_inb = 147;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 148;
address_inb = 149;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 150;
address_inb = 151;
data_ina = 16'h2;
data_inb = 16'h0;
#10;
address_ina = 152;
address_inb = 153;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 154;
address_inb = 155;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 156;
address_inb = 157;
data_ina = 16'h0;
data_inb = 16'hfffe;
#10;
address_ina = 158;
address_inb = 159;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 160;
address_inb = 161;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 162;
address_inb = 163;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 164;
address_inb = 165;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 166;
address_inb = 167;
data_ina = 16'h2;
data_inb = 16'h0;
#10;
address_ina = 168;
address_inb = 169;
data_ina = 16'hffff;
data_inb = 16'h2;
#10;
address_ina = 170;
address_inb = 171;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 172;
address_inb = 173;
data_ina = 16'hffff;
data_inb = 16'hfffe;
#10;
address_ina = 174;
address_inb = 175;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 176;
address_inb = 177;
data_ina = 16'h2;
data_inb = 16'h2;
#10;
address_ina = 178;
address_inb = 179;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 180;
address_inb = 181;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 182;
address_inb = 183;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 184;
address_inb = 185;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 186;
address_inb = 187;
data_ina = 16'h3;
data_inb = 16'h0;
#10;
address_ina = 188;
address_inb = 189;
data_ina = 16'hfffe;
data_inb = 16'h3;
#10;
address_ina = 190;
address_inb = 191;
data_ina = 16'h0;
data_inb = 16'h2;
#10;
address_ina = 192;
address_inb = 193;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 194;
address_inb = 195;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 196;
address_inb = 197;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 198;
address_inb = 199;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 200;
address_inb = 201;
data_ina = 16'hfffe;
data_inb = 16'h1;
#10;
address_ina = 202;
address_inb = 203;
data_ina = 16'h0;
data_inb = 16'h2;
#10;
address_ina = 204;
address_inb = 205;
data_ina = 16'h0;
data_inb = 16'hfffe;
#10;
address_ina = 206;
address_inb = 207;
data_ina = 16'h2;
data_inb = 16'h0;
#10;
address_ina = 208;
address_inb = 209;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 210;
address_inb = 211;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 212;
address_inb = 213;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 214;
address_inb = 215;
data_ina = 16'hfffd;
data_inb = 16'hffff;
#10;
address_ina = 216;
address_inb = 217;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 218;
address_inb = 219;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 220;
address_inb = 221;
data_ina = 16'hfffe;
data_inb = 16'h0;
#10;
address_ina = 222;
address_inb = 223;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 224;
address_inb = 225;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 226;
address_inb = 227;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 228;
address_inb = 229;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 230;
address_inb = 231;
data_ina = 16'h2;
data_inb = 16'h1;
#10;
address_ina = 232;
address_inb = 233;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 234;
address_inb = 235;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 236;
address_inb = 237;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 238;
address_inb = 239;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 240;
address_inb = 241;
data_ina = 16'h0;
data_inb = 16'hfffe;
#10;
address_ina = 242;
address_inb = 243;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 244;
address_inb = 245;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 246;
address_inb = 247;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 248;
address_inb = 249;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 250;
address_inb = 251;
data_ina = 16'h2;
data_inb = 16'h3;
#10;
address_ina = 252;
address_inb = 253;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 254;
address_inb = 255;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
        wait(init_done);
        #30
        we = 0;
        // Start processing
         
		  #38000

        start = 0;



//        wait (wr_req);
//		  wait (!wr_req);
//		   rd_req = 1;
		  wait(done);
		  #20000
rd_req = 1;
        #70 
		  start = 1;
		 #80 
wait(rd_empty)
rd_req = 0;

$display("Finished the NTT test Number %d",test_num);
////Begin test number #47//////////////
rst = 1;

//#1000
start = 1;
mode = 0; //NTT 0 // INTT 1

// Reset for a few clock cycles

#1000

rst = 0;
test_num = test_num + 1;
#1000
we = 1;
address_ina = 0;
address_inb = 1;
data_ina = 16'h1;
data_inb = 16'hfffe;
#10;
address_ina = 2;
address_inb = 3;
data_ina = 16'h2;
data_inb = 16'hffff;
#10;
address_ina = 4;
address_inb = 5;
data_ina = 16'hfffe;
data_inb = 16'hffff;
#10;
address_ina = 6;
address_inb = 7;
data_ina = 16'h2;
data_inb = 16'h0;
#10;
address_ina = 8;
address_inb = 9;
data_ina = 16'hfffe;
data_inb = 16'h0;
#10;
address_ina = 10;
address_inb = 11;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 12;
address_inb = 13;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 14;
address_inb = 15;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 16;
address_inb = 17;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 18;
address_inb = 19;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 20;
address_inb = 21;
data_ina = 16'hfffe;
data_inb = 16'h1;
#10;
address_ina = 22;
address_inb = 23;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 24;
address_inb = 25;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 26;
address_inb = 27;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 28;
address_inb = 29;
data_ina = 16'hffff;
data_inb = 16'hfffe;
#10;
address_ina = 30;
address_inb = 31;
data_ina = 16'h2;
data_inb = 16'hfffe;
#10;
address_ina = 32;
address_inb = 33;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 34;
address_inb = 35;
data_ina = 16'h2;
data_inb = 16'h0;
#10;
address_ina = 36;
address_inb = 37;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 38;
address_inb = 39;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 40;
address_inb = 41;
data_ina = 16'h2;
data_inb = 16'h3;
#10;
address_ina = 42;
address_inb = 43;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 44;
address_inb = 45;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 46;
address_inb = 47;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 48;
address_inb = 49;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 50;
address_inb = 51;
data_ina = 16'h1;
data_inb = 16'hfffe;
#10;
address_ina = 52;
address_inb = 53;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 54;
address_inb = 55;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 56;
address_inb = 57;
data_ina = 16'hfffe;
data_inb = 16'hffff;
#10;
address_ina = 58;
address_inb = 59;
data_ina = 16'hffff;
data_inb = 16'h2;
#10;
address_ina = 60;
address_inb = 61;
data_ina = 16'hfffe;
data_inb = 16'h0;
#10;
address_ina = 62;
address_inb = 63;
data_ina = 16'hffff;
data_inb = 16'h2;
#10;
address_ina = 64;
address_inb = 65;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 66;
address_inb = 67;
data_ina = 16'h2;
data_inb = 16'h0;
#10;
address_ina = 68;
address_inb = 69;
data_ina = 16'h0;
data_inb = 16'hfffe;
#10;
address_ina = 70;
address_inb = 71;
data_ina = 16'h1;
data_inb = 16'h2;
#10;
address_ina = 72;
address_inb = 73;
data_ina = 16'hfffd;
data_inb = 16'h0;
#10;
address_ina = 74;
address_inb = 75;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 76;
address_inb = 77;
data_ina = 16'hfffe;
data_inb = 16'h0;
#10;
address_ina = 78;
address_inb = 79;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 80;
address_inb = 81;
data_ina = 16'hfffe;
data_inb = 16'hffff;
#10;
address_ina = 82;
address_inb = 83;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 84;
address_inb = 85;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 86;
address_inb = 87;
data_ina = 16'hfffe;
data_inb = 16'h2;
#10;
address_ina = 88;
address_inb = 89;
data_ina = 16'hfffd;
data_inb = 16'h1;
#10;
address_ina = 90;
address_inb = 91;
data_ina = 16'h0;
data_inb = 16'hfffe;
#10;
address_ina = 92;
address_inb = 93;
data_ina = 16'h0;
data_inb = 16'h3;
#10;
address_ina = 94;
address_inb = 95;
data_ina = 16'hfffe;
data_inb = 16'h2;
#10;
address_ina = 96;
address_inb = 97;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 98;
address_inb = 99;
data_ina = 16'hfffe;
data_inb = 16'hfffe;
#10;
address_ina = 100;
address_inb = 101;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 102;
address_inb = 103;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 104;
address_inb = 105;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 106;
address_inb = 107;
data_ina = 16'h0;
data_inb = 16'h3;
#10;
address_ina = 108;
address_inb = 109;
data_ina = 16'h0;
data_inb = 16'hfffe;
#10;
address_ina = 110;
address_inb = 111;
data_ina = 16'h1;
data_inb = 16'hfffe;
#10;
address_ina = 112;
address_inb = 113;
data_ina = 16'h2;
data_inb = 16'h0;
#10;
address_ina = 114;
address_inb = 115;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 116;
address_inb = 117;
data_ina = 16'h0;
data_inb = 16'h3;
#10;
address_ina = 118;
address_inb = 119;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 120;
address_inb = 121;
data_ina = 16'hffff;
data_inb = 16'hfffe;
#10;
address_ina = 122;
address_inb = 123;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 124;
address_inb = 125;
data_ina = 16'hfffe;
data_inb = 16'hffff;
#10;
address_ina = 126;
address_inb = 127;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 128;
address_inb = 129;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 130;
address_inb = 131;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 132;
address_inb = 133;
data_ina = 16'h1;
data_inb = 16'hfffe;
#10;
address_ina = 134;
address_inb = 135;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 136;
address_inb = 137;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 138;
address_inb = 139;
data_ina = 16'hfffe;
data_inb = 16'h0;
#10;
address_ina = 140;
address_inb = 141;
data_ina = 16'h1;
data_inb = 16'hfffe;
#10;
address_ina = 142;
address_inb = 143;
data_ina = 16'hffff;
data_inb = 16'h2;
#10;
address_ina = 144;
address_inb = 145;
data_ina = 16'h2;
data_inb = 16'h0;
#10;
address_ina = 146;
address_inb = 147;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 148;
address_inb = 149;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 150;
address_inb = 151;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 152;
address_inb = 153;
data_ina = 16'hffff;
data_inb = 16'h2;
#10;
address_ina = 154;
address_inb = 155;
data_ina = 16'h0;
data_inb = 16'h2;
#10;
address_ina = 156;
address_inb = 157;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 158;
address_inb = 159;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 160;
address_inb = 161;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 162;
address_inb = 163;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 164;
address_inb = 165;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 166;
address_inb = 167;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 168;
address_inb = 169;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 170;
address_inb = 171;
data_ina = 16'h2;
data_inb = 16'h0;
#10;
address_ina = 172;
address_inb = 173;
data_ina = 16'hffff;
data_inb = 16'hfffe;
#10;
address_ina = 174;
address_inb = 175;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 176;
address_inb = 177;
data_ina = 16'h2;
data_inb = 16'h0;
#10;
address_ina = 178;
address_inb = 179;
data_ina = 16'h2;
data_inb = 16'h1;
#10;
address_ina = 180;
address_inb = 181;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 182;
address_inb = 183;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 184;
address_inb = 185;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 186;
address_inb = 187;
data_ina = 16'hffff;
data_inb = 16'h2;
#10;
address_ina = 188;
address_inb = 189;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 190;
address_inb = 191;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 192;
address_inb = 193;
data_ina = 16'h0;
data_inb = 16'hfffe;
#10;
address_ina = 194;
address_inb = 195;
data_ina = 16'h1;
data_inb = 16'h2;
#10;
address_ina = 196;
address_inb = 197;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 198;
address_inb = 199;
data_ina = 16'hffff;
data_inb = 16'hfffe;
#10;
address_ina = 200;
address_inb = 201;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 202;
address_inb = 203;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 204;
address_inb = 205;
data_ina = 16'h0;
data_inb = 16'h3;
#10;
address_ina = 206;
address_inb = 207;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 208;
address_inb = 209;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 210;
address_inb = 211;
data_ina = 16'h2;
data_inb = 16'h2;
#10;
address_ina = 212;
address_inb = 213;
data_ina = 16'h2;
data_inb = 16'h1;
#10;
address_ina = 214;
address_inb = 215;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 216;
address_inb = 217;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 218;
address_inb = 219;
data_ina = 16'hfffe;
data_inb = 16'h0;
#10;
address_ina = 220;
address_inb = 221;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 222;
address_inb = 223;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 224;
address_inb = 225;
data_ina = 16'h2;
data_inb = 16'h0;
#10;
address_ina = 226;
address_inb = 227;
data_ina = 16'h3;
data_inb = 16'h0;
#10;
address_ina = 228;
address_inb = 229;
data_ina = 16'hfffe;
data_inb = 16'h1;
#10;
address_ina = 230;
address_inb = 231;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 232;
address_inb = 233;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 234;
address_inb = 235;
data_ina = 16'hffff;
data_inb = 16'hfffe;
#10;
address_ina = 236;
address_inb = 237;
data_ina = 16'hffff;
data_inb = 16'hfffe;
#10;
address_ina = 238;
address_inb = 239;
data_ina = 16'hffff;
data_inb = 16'hfffe;
#10;
address_ina = 240;
address_inb = 241;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 242;
address_inb = 243;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 244;
address_inb = 245;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 246;
address_inb = 247;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 248;
address_inb = 249;
data_ina = 16'hfffe;
data_inb = 16'h2;
#10;
address_ina = 250;
address_inb = 251;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 252;
address_inb = 253;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 254;
address_inb = 255;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
        wait(init_done);
        #30
        we = 0;
        // Start processing
         
		  #38000

        start = 0;



//        wait (wr_req);
//		  wait (!wr_req);
//		   rd_req = 1;
		  wait(done);
		  #20000
rd_req = 1;
        #70 
		  start = 1;
		 #80 
wait(rd_empty)
rd_req = 0;

$display("Finished the NTT test Number %d",test_num);
////Begin test number #48//////////////
rst = 1;

//#1000
start = 1;
mode = 1; //NTT 0 // INTT 1

// Reset for a few clock cycles

#1000

rst = 0;
test_num = test_num + 1;
#1000
we = 1;
address_ina = 0;
address_inb = 1;
data_ina = 16'hf9e0;
data_inb = 16'hfa0e;
#10;
address_ina = 2;
address_inb = 3;
data_ina = 16'h43;
data_inb = 16'hfb61;
#10;
address_ina = 4;
address_inb = 5;
data_ina = 16'h2f7;
data_inb = 16'hff7d;
#10;
address_ina = 6;
address_inb = 7;
data_ina = 16'h5c6;
data_inb = 16'h29d;
#10;
address_ina = 8;
address_inb = 9;
data_ina = 16'hfc52;
data_inb = 16'hff76;
#10;
address_ina = 10;
address_inb = 11;
data_ina = 16'h4fa;
data_inb = 16'h2ef;
#10;
address_ina = 12;
address_inb = 13;
data_ina = 16'h555;
data_inb = 16'h4fd;
#10;
address_ina = 14;
address_inb = 15;
data_ina = 16'hfdc3;
data_inb = 16'hfec1;
#10;
address_ina = 16;
address_inb = 17;
data_ina = 16'h54d;
data_inb = 16'h5d0;
#10;
address_ina = 18;
address_inb = 19;
data_ina = 16'h454;
data_inb = 16'hff6d;
#10;
address_ina = 20;
address_inb = 21;
data_ina = 16'hfb53;
data_inb = 16'hffd9;
#10;
address_ina = 22;
address_inb = 23;
data_ina = 16'he9;
data_inb = 16'hfce4;
#10;
address_ina = 24;
address_inb = 25;
data_ina = 16'hfb46;
data_inb = 16'h65d;
#10;
address_ina = 26;
address_inb = 27;
data_ina = 16'hffcf;
data_inb = 16'hfe85;
#10;
address_ina = 28;
address_inb = 29;
data_ina = 16'h174;
data_inb = 16'h15a;
#10;
address_ina = 30;
address_inb = 31;
data_ina = 16'h129;
data_inb = 16'hfaa8;
#10;
address_ina = 32;
address_inb = 33;
data_ina = 16'hfe3e;
data_inb = 16'h72;
#10;
address_ina = 34;
address_inb = 35;
data_ina = 16'hfb02;
data_inb = 16'h3e3;
#10;
address_ina = 36;
address_inb = 37;
data_ina = 16'h30e;
data_inb = 16'h10a;
#10;
address_ina = 38;
address_inb = 39;
data_ina = 16'hfbcc;
data_inb = 16'hfdc1;
#10;
address_ina = 40;
address_inb = 41;
data_ina = 16'hff11;
data_inb = 16'h5ad;
#10;
address_ina = 42;
address_inb = 43;
data_ina = 16'h676;
data_inb = 16'hfb16;
#10;
address_ina = 44;
address_inb = 45;
data_ina = 16'haa;
data_inb = 16'hfed1;
#10;
address_ina = 46;
address_inb = 47;
data_ina = 16'hfcdc;
data_inb = 16'hfbc6;
#10;
address_ina = 48;
address_inb = 49;
data_ina = 16'h43f;
data_inb = 16'hfb1f;
#10;
address_ina = 50;
address_inb = 51;
data_ina = 16'h193;
data_inb = 16'h5d7;
#10;
address_ina = 52;
address_inb = 53;
data_ina = 16'hfd89;
data_inb = 16'h294;
#10;
address_ina = 54;
address_inb = 55;
data_ina = 16'h577;
data_inb = 16'hfbc5;
#10;
address_ina = 56;
address_inb = 57;
data_ina = 16'hc9;
data_inb = 16'hfd6b;
#10;
address_ina = 58;
address_inb = 59;
data_ina = 16'h1f0;
data_inb = 16'h472;
#10;
address_ina = 60;
address_inb = 61;
data_ina = 16'h5c9;
data_inb = 16'h5d9;
#10;
address_ina = 62;
address_inb = 63;
data_ina = 16'hfcb0;
data_inb = 16'h3cf;
#10;
address_ina = 64;
address_inb = 65;
data_ina = 16'hfe61;
data_inb = 16'hfef8;
#10;
address_ina = 66;
address_inb = 67;
data_ina = 16'h176;
data_inb = 16'hfbff;
#10;
address_ina = 68;
address_inb = 69;
data_ina = 16'h1df;
data_inb = 16'h4b2;
#10;
address_ina = 70;
address_inb = 71;
data_ina = 16'hfacd;
data_inb = 16'h1e8;
#10;
address_ina = 72;
address_inb = 73;
data_ina = 16'h5d2;
data_inb = 16'h2d6;
#10;
address_ina = 74;
address_inb = 75;
data_ina = 16'h144;
data_inb = 16'hfcd8;
#10;
address_ina = 76;
address_inb = 77;
data_ina = 16'h8e;
data_inb = 16'hf9d4;
#10;
address_ina = 78;
address_inb = 79;
data_ina = 16'hfb7d;
data_inb = 16'hf9ed;
#10;
address_ina = 80;
address_inb = 81;
data_ina = 16'hfd10;
data_inb = 16'hfc67;
#10;
address_ina = 82;
address_inb = 83;
data_ina = 16'hfe64;
data_inb = 16'hffa2;
#10;
address_ina = 84;
address_inb = 85;
data_ina = 16'h52d;
data_inb = 16'hea;
#10;
address_ina = 86;
address_inb = 87;
data_ina = 16'h37c;
data_inb = 16'hfebe;
#10;
address_ina = 88;
address_inb = 89;
data_ina = 16'h36a;
data_inb = 16'hfd33;
#10;
address_ina = 90;
address_inb = 91;
data_ina = 16'h158;
data_inb = 16'h30;
#10;
address_ina = 92;
address_inb = 93;
data_ina = 16'h618;
data_inb = 16'hfbb3;
#10;
address_ina = 94;
address_inb = 95;
data_ina = 16'hfdd2;
data_inb = 16'hfd1d;
#10;
address_ina = 96;
address_inb = 97;
data_ina = 16'hfc9a;
data_inb = 16'hfdec;
#10;
address_ina = 98;
address_inb = 99;
data_ina = 16'hfdd4;
data_inb = 16'hfe21;
#10;
address_ina = 100;
address_inb = 101;
data_ina = 16'h643;
data_inb = 16'hfbc5;
#10;
address_ina = 102;
address_inb = 103;
data_ina = 16'hfce2;
data_inb = 16'h206;
#10;
address_ina = 104;
address_inb = 105;
data_ina = 16'hfe00;
data_inb = 16'h2db;
#10;
address_ina = 106;
address_inb = 107;
data_ina = 16'h58;
data_inb = 16'h2e6;
#10;
address_ina = 108;
address_inb = 109;
data_ina = 16'hfb7c;
data_inb = 16'hfd14;
#10;
address_ina = 110;
address_inb = 111;
data_ina = 16'h430;
data_inb = 16'hfe9b;
#10;
address_ina = 112;
address_inb = 113;
data_ina = 16'hfa5a;
data_inb = 16'h31e;
#10;
address_ina = 114;
address_inb = 115;
data_ina = 16'h599;
data_inb = 16'h5a5;
#10;
address_ina = 116;
address_inb = 117;
data_ina = 16'h30b;
data_inb = 16'hfa56;
#10;
address_ina = 118;
address_inb = 119;
data_ina = 16'h573;
data_inb = 16'hfc3e;
#10;
address_ina = 120;
address_inb = 121;
data_ina = 16'hff62;
data_inb = 16'hfc69;
#10;
address_ina = 122;
address_inb = 123;
data_ina = 16'hf99d;
data_inb = 16'h654;
#10;
address_ina = 124;
address_inb = 125;
data_ina = 16'h3a9;
data_inb = 16'h322;
#10;
address_ina = 126;
address_inb = 127;
data_ina = 16'hfd6a;
data_inb = 16'hfa7c;
#10;
address_ina = 128;
address_inb = 129;
data_ina = 16'hfcc3;
data_inb = 16'hfe7f;
#10;
address_ina = 130;
address_inb = 131;
data_ina = 16'h403;
data_inb = 16'hfbde;
#10;
address_ina = 132;
address_inb = 133;
data_ina = 16'hfa89;
data_inb = 16'hfe2e;
#10;
address_ina = 134;
address_inb = 135;
data_ina = 16'hfe2d;
data_inb = 16'hfb0c;
#10;
address_ina = 136;
address_inb = 137;
data_ina = 16'h21e;
data_inb = 16'h58d;
#10;
address_ina = 138;
address_inb = 139;
data_ina = 16'h18d;
data_inb = 16'hfae9;
#10;
address_ina = 140;
address_inb = 141;
data_ina = 16'h7;
data_inb = 16'hfef8;
#10;
address_ina = 142;
address_inb = 143;
data_ina = 16'hfe1d;
data_inb = 16'h30f;
#10;
address_ina = 144;
address_inb = 145;
data_ina = 16'h11b;
data_inb = 16'h486;
#10;
address_ina = 146;
address_inb = 147;
data_ina = 16'hfcb6;
data_inb = 16'h43;
#10;
address_ina = 148;
address_inb = 149;
data_ina = 16'hfb43;
data_inb = 16'h243;
#10;
address_ina = 150;
address_inb = 151;
data_ina = 16'h84;
data_inb = 16'h555;
#10;
address_ina = 152;
address_inb = 153;
data_ina = 16'h372;
data_inb = 16'h222;
#10;
address_ina = 154;
address_inb = 155;
data_ina = 16'hfcd6;
data_inb = 16'hfe8b;
#10;
address_ina = 156;
address_inb = 157;
data_ina = 16'h5ef;
data_inb = 16'hfe51;
#10;
address_ina = 158;
address_inb = 159;
data_ina = 16'hfc24;
data_inb = 16'h1e;
#10;
address_ina = 160;
address_inb = 161;
data_ina = 16'h60e;
data_inb = 16'hff;
#10;
address_ina = 162;
address_inb = 163;
data_ina = 16'hfe1d;
data_inb = 16'h480;
#10;
address_ina = 164;
address_inb = 165;
data_ina = 16'hfc19;
data_inb = 16'hfcb5;
#10;
address_ina = 166;
address_inb = 167;
data_ina = 16'h221;
data_inb = 16'h43f;
#10;
address_ina = 168;
address_inb = 169;
data_ina = 16'hfccf;
data_inb = 16'hfc47;
#10;
address_ina = 170;
address_inb = 171;
data_ina = 16'h1fe;
data_inb = 16'hf9ff;
#10;
address_ina = 172;
address_inb = 173;
data_ina = 16'hfe38;
data_inb = 16'h5da;
#10;
address_ina = 174;
address_inb = 175;
data_ina = 16'h132;
data_inb = 16'hfdac;
#10;
address_ina = 176;
address_inb = 177;
data_ina = 16'h673;
data_inb = 16'hf9ba;
#10;
address_ina = 178;
address_inb = 179;
data_ina = 16'hfd19;
data_inb = 16'hfe72;
#10;
address_ina = 180;
address_inb = 181;
data_ina = 16'hfec3;
data_inb = 16'hfde6;
#10;
address_ina = 182;
address_inb = 183;
data_ina = 16'hfcd6;
data_inb = 16'h390;
#10;
address_ina = 184;
address_inb = 185;
data_ina = 16'hfd26;
data_inb = 16'h372;
#10;
address_ina = 186;
address_inb = 187;
data_ina = 16'h50b;
data_inb = 16'h248;
#10;
address_ina = 188;
address_inb = 189;
data_ina = 16'h4f4;
data_inb = 16'h88;
#10;
address_ina = 190;
address_inb = 191;
data_ina = 16'h3ed;
data_inb = 16'h1b1;
#10;
address_ina = 192;
address_inb = 193;
data_ina = 16'h5b8;
data_inb = 16'h81;
#10;
address_ina = 194;
address_inb = 195;
data_ina = 16'hfc53;
data_inb = 16'h546;
#10;
address_ina = 196;
address_inb = 197;
data_ina = 16'h3c9;
data_inb = 16'h3e9;
#10;
address_ina = 198;
address_inb = 199;
data_ina = 16'hf994;
data_inb = 16'h4da;
#10;
address_ina = 200;
address_inb = 201;
data_ina = 16'hfa89;
data_inb = 16'hfe0f;
#10;
address_ina = 202;
address_inb = 203;
data_ina = 16'h4a5;
data_inb = 16'hfb53;
#10;
address_ina = 204;
address_inb = 205;
data_ina = 16'h1be;
data_inb = 16'hff81;
#10;
address_ina = 206;
address_inb = 207;
data_ina = 16'hfa35;
data_inb = 16'h314;
#10;
address_ina = 208;
address_inb = 209;
data_ina = 16'hfdec;
data_inb = 16'h343;
#10;
address_ina = 210;
address_inb = 211;
data_ina = 16'h552;
data_inb = 16'h25;
#10;
address_ina = 212;
address_inb = 213;
data_ina = 16'h51d;
data_inb = 16'hff40;
#10;
address_ina = 214;
address_inb = 215;
data_ina = 16'h551;
data_inb = 16'hfc2a;
#10;
address_ina = 216;
address_inb = 217;
data_ina = 16'h5d3;
data_inb = 16'h5be;
#10;
address_ina = 218;
address_inb = 219;
data_ina = 16'h50a;
data_inb = 16'hfa32;
#10;
address_ina = 220;
address_inb = 221;
data_ina = 16'hb3;
data_inb = 16'h158;
#10;
address_ina = 222;
address_inb = 223;
data_ina = 16'hfcc0;
data_inb = 16'hfb26;
#10;
address_ina = 224;
address_inb = 225;
data_ina = 16'h5a0;
data_inb = 16'hfbaf;
#10;
address_ina = 226;
address_inb = 227;
data_ina = 16'hfdeb;
data_inb = 16'hf9dc;
#10;
address_ina = 228;
address_inb = 229;
data_ina = 16'hfadd;
data_inb = 16'hff33;
#10;
address_ina = 230;
address_inb = 231;
data_ina = 16'hfcaa;
data_inb = 16'hff13;
#10;
address_ina = 232;
address_inb = 233;
data_ina = 16'h335;
data_inb = 16'h3e3;
#10;
address_ina = 234;
address_inb = 235;
data_ina = 16'hf9e4;
data_inb = 16'hfe1e;
#10;
address_ina = 236;
address_inb = 237;
data_ina = 16'h322;
data_inb = 16'h5d1;
#10;
address_ina = 238;
address_inb = 239;
data_ina = 16'h3f7;
data_inb = 16'hfb19;
#10;
address_ina = 240;
address_inb = 241;
data_ina = 16'hfd19;
data_inb = 16'hfc38;
#10;
address_ina = 242;
address_inb = 243;
data_ina = 16'h48c;
data_inb = 16'h45d;
#10;
address_ina = 244;
address_inb = 245;
data_ina = 16'hfb1a;
data_inb = 16'h4d6;
#10;
address_ina = 246;
address_inb = 247;
data_ina = 16'h101;
data_inb = 16'hfae1;
#10;
address_ina = 248;
address_inb = 249;
data_ina = 16'hfc18;
data_inb = 16'h369;
#10;
address_ina = 250;
address_inb = 251;
data_ina = 16'h1b0;
data_inb = 16'h185;
#10;
address_ina = 252;
address_inb = 253;
data_ina = 16'h28f;
data_inb = 16'hfae9;
#10;
address_ina = 254;
address_inb = 255;
data_ina = 16'hfbc0;
data_inb = 16'h2b4;
#10;
        wait(init_done);
        #30
        we = 0;
        // Start processing
         
		  #38000

        start = 0;



//        wait (wr_req);
//		  wait (!wr_req);
//		   rd_req = 1;
		  wait(done);
		  #20000
rd_req = 1;
        #70 
		  start = 1;
		 #80 
wait(rd_empty)
rd_req = 0;

$display("Finished the NTT test Number %d",test_num);
////Begin test number #49//////////////
rst = 1;

//#1000
start = 1;
mode = 1; //NTT 0 // INTT 1

// Reset for a few clock cycles

#1000

rst = 0;
test_num = test_num + 1;
#1000
we = 1;
address_ina = 0;
address_inb = 1;
data_ina = 16'h582;
data_inb = 16'hfa79;
#10;
address_ina = 2;
address_inb = 3;
data_ina = 16'hfd8d;
data_inb = 16'hfad4;
#10;
address_ina = 4;
address_inb = 5;
data_ina = 16'h1b8;
data_inb = 16'hff;
#10;
address_ina = 6;
address_inb = 7;
data_ina = 16'hfa3c;
data_inb = 16'h3d2;
#10;
address_ina = 8;
address_inb = 9;
data_ina = 16'hff83;
data_inb = 16'h460;
#10;
address_ina = 10;
address_inb = 11;
data_ina = 16'hfdb0;
data_inb = 16'h5a3;
#10;
address_ina = 12;
address_inb = 13;
data_ina = 16'h3b2;
data_inb = 16'hfdea;
#10;
address_ina = 14;
address_inb = 15;
data_ina = 16'hfb27;
data_inb = 16'h107;
#10;
address_ina = 16;
address_inb = 17;
data_ina = 16'hffbb;
data_inb = 16'h511;
#10;
address_ina = 18;
address_inb = 19;
data_ina = 16'h2b9;
data_inb = 16'hfcda;
#10;
address_ina = 20;
address_inb = 21;
data_ina = 16'hff35;
data_inb = 16'hfa9e;
#10;
address_ina = 22;
address_inb = 23;
data_ina = 16'hfc43;
data_inb = 16'hfd32;
#10;
address_ina = 24;
address_inb = 25;
data_ina = 16'h1d4;
data_inb = 16'hc6;
#10;
address_ina = 26;
address_inb = 27;
data_ina = 16'hfe27;
data_inb = 16'h557;
#10;
address_ina = 28;
address_inb = 29;
data_ina = 16'hfb2c;
data_inb = 16'h318;
#10;
address_ina = 30;
address_inb = 31;
data_ina = 16'h1f8;
data_inb = 16'hfe2b;
#10;
address_ina = 32;
address_inb = 33;
data_ina = 16'h633;
data_inb = 16'hfbcd;
#10;
address_ina = 34;
address_inb = 35;
data_ina = 16'hf9f8;
data_inb = 16'h41f;
#10;
address_ina = 36;
address_inb = 37;
data_ina = 16'hfe9d;
data_inb = 16'h35c;
#10;
address_ina = 38;
address_inb = 39;
data_ina = 16'h1c7;
data_inb = 16'h35f;
#10;
address_ina = 40;
address_inb = 41;
data_ina = 16'h637;
data_inb = 16'h57;
#10;
address_ina = 42;
address_inb = 43;
data_ina = 16'h313;
data_inb = 16'hfc2d;
#10;
address_ina = 44;
address_inb = 45;
data_ina = 16'ha2;
data_inb = 16'h65c;
#10;
address_ina = 46;
address_inb = 47;
data_ina = 16'h326;
data_inb = 16'hf9c0;
#10;
address_ina = 48;
address_inb = 49;
data_ina = 16'h4e4;
data_inb = 16'h4fc;
#10;
address_ina = 50;
address_inb = 51;
data_ina = 16'hfc01;
data_inb = 16'hfaa5;
#10;
address_ina = 52;
address_inb = 53;
data_ina = 16'h62d;
data_inb = 16'hfda0;
#10;
address_ina = 54;
address_inb = 55;
data_ina = 16'h662;
data_inb = 16'h44d;
#10;
address_ina = 56;
address_inb = 57;
data_ina = 16'hf9d0;
data_inb = 16'hdb;
#10;
address_ina = 58;
address_inb = 59;
data_ina = 16'hf984;
data_inb = 16'h37f;
#10;
address_ina = 60;
address_inb = 61;
data_ina = 16'hf9cf;
data_inb = 16'h2b4;
#10;
address_ina = 62;
address_inb = 63;
data_ina = 16'hfd59;
data_inb = 16'hfe0f;
#10;
address_ina = 64;
address_inb = 65;
data_ina = 16'h62b;
data_inb = 16'h4ee;
#10;
address_ina = 66;
address_inb = 67;
data_ina = 16'hfc5e;
data_inb = 16'h504;
#10;
address_ina = 68;
address_inb = 69;
data_ina = 16'hffab;
data_inb = 16'hff08;
#10;
address_ina = 70;
address_inb = 71;
data_ina = 16'h23c;
data_inb = 16'hfc1f;
#10;
address_ina = 72;
address_inb = 73;
data_ina = 16'hfe6c;
data_inb = 16'h5dc;
#10;
address_ina = 74;
address_inb = 75;
data_ina = 16'hfea1;
data_inb = 16'h5d3;
#10;
address_ina = 76;
address_inb = 77;
data_ina = 16'hc8;
data_inb = 16'hf9df;
#10;
address_ina = 78;
address_inb = 79;
data_ina = 16'h40d;
data_inb = 16'h512;
#10;
address_ina = 80;
address_inb = 81;
data_ina = 16'h616;
data_inb = 16'hfe57;
#10;
address_ina = 82;
address_inb = 83;
data_ina = 16'hfc44;
data_inb = 16'h95;
#10;
address_ina = 84;
address_inb = 85;
data_ina = 16'hfc90;
data_inb = 16'hfb66;
#10;
address_ina = 86;
address_inb = 87;
data_ina = 16'h35d;
data_inb = 16'h45b;
#10;
address_ina = 88;
address_inb = 89;
data_ina = 16'hfdac;
data_inb = 16'h2bb;
#10;
address_ina = 90;
address_inb = 91;
data_ina = 16'h90;
data_inb = 16'h138;
#10;
address_ina = 92;
address_inb = 93;
data_ina = 16'hfbc8;
data_inb = 16'h5c0;
#10;
address_ina = 94;
address_inb = 95;
data_ina = 16'h58;
data_inb = 16'hfe0b;
#10;
address_ina = 96;
address_inb = 97;
data_ina = 16'hfe8b;
data_inb = 16'hffe0;
#10;
address_ina = 98;
address_inb = 99;
data_ina = 16'hffd8;
data_inb = 16'hfdaf;
#10;
address_ina = 100;
address_inb = 101;
data_ina = 16'h5e2;
data_inb = 16'hfd95;
#10;
address_ina = 102;
address_inb = 103;
data_ina = 16'hfc71;
data_inb = 16'hfdb9;
#10;
address_ina = 104;
address_inb = 105;
data_ina = 16'h5a7;
data_inb = 16'hffea;
#10;
address_ina = 106;
address_inb = 107;
data_ina = 16'h3e7;
data_inb = 16'h2a8;
#10;
address_ina = 108;
address_inb = 109;
data_ina = 16'h51c;
data_inb = 16'hfc74;
#10;
address_ina = 110;
address_inb = 111;
data_ina = 16'hfcc7;
data_inb = 16'h4dd;
#10;
address_ina = 112;
address_inb = 113;
data_ina = 16'h5ad;
data_inb = 16'hfc3c;
#10;
address_ina = 114;
address_inb = 115;
data_ina = 16'hfd9d;
data_inb = 16'h52c;
#10;
address_ina = 116;
address_inb = 117;
data_ina = 16'h16b;
data_inb = 16'hffcb;
#10;
address_ina = 118;
address_inb = 119;
data_ina = 16'hfcfc;
data_inb = 16'hfb6e;
#10;
address_ina = 120;
address_inb = 121;
data_ina = 16'hfd55;
data_inb = 16'hfa58;
#10;
address_ina = 122;
address_inb = 123;
data_ina = 16'hfb29;
data_inb = 16'h35a;
#10;
address_ina = 124;
address_inb = 125;
data_ina = 16'h474;
data_inb = 16'h2e8;
#10;
address_ina = 126;
address_inb = 127;
data_ina = 16'h298;
data_inb = 16'hfcc8;
#10;
address_ina = 128;
address_inb = 129;
data_ina = 16'hfc71;
data_inb = 16'hfd66;
#10;
address_ina = 130;
address_inb = 131;
data_ina = 16'h4e3;
data_inb = 16'hfacb;
#10;
address_ina = 132;
address_inb = 133;
data_ina = 16'hf9ae;
data_inb = 16'h5b2;
#10;
address_ina = 134;
address_inb = 135;
data_ina = 16'h49d;
data_inb = 16'h457;
#10;
address_ina = 136;
address_inb = 137;
data_ina = 16'hffeb;
data_inb = 16'h328;
#10;
address_ina = 138;
address_inb = 139;
data_ina = 16'h3ec;
data_inb = 16'hfd4e;
#10;
address_ina = 140;
address_inb = 141;
data_ina = 16'h418;
data_inb = 16'hfc63;
#10;
address_ina = 142;
address_inb = 143;
data_ina = 16'h1a8;
data_inb = 16'h44a;
#10;
address_ina = 144;
address_inb = 145;
data_ina = 16'hff95;
data_inb = 16'hfc62;
#10;
address_ina = 146;
address_inb = 147;
data_ina = 16'h42f;
data_inb = 16'h624;
#10;
address_ina = 148;
address_inb = 149;
data_ina = 16'hfdfe;
data_inb = 16'h388;
#10;
address_ina = 150;
address_inb = 151;
data_ina = 16'hfc7d;
data_inb = 16'h64e;
#10;
address_ina = 152;
address_inb = 153;
data_ina = 16'hfe3a;
data_inb = 16'h1ce;
#10;
address_ina = 154;
address_inb = 155;
data_ina = 16'hfe94;
data_inb = 16'hfc34;
#10;
address_ina = 156;
address_inb = 157;
data_ina = 16'hff07;
data_inb = 16'hfcb1;
#10;
address_ina = 158;
address_inb = 159;
data_ina = 16'hfc46;
data_inb = 16'h157;
#10;
address_ina = 160;
address_inb = 161;
data_ina = 16'h1e6;
data_inb = 16'hfdb3;
#10;
address_ina = 162;
address_inb = 163;
data_ina = 16'hfda7;
data_inb = 16'hfb81;
#10;
address_ina = 164;
address_inb = 165;
data_ina = 16'hf9d4;
data_inb = 16'hfb88;
#10;
address_ina = 166;
address_inb = 167;
data_ina = 16'hfe79;
data_inb = 16'h488;
#10;
address_ina = 168;
address_inb = 169;
data_ina = 16'hfebc;
data_inb = 16'hfeb1;
#10;
address_ina = 170;
address_inb = 171;
data_ina = 16'hfbe4;
data_inb = 16'hfe78;
#10;
address_ina = 172;
address_inb = 173;
data_ina = 16'h67d;
data_inb = 16'h3ed;
#10;
address_ina = 174;
address_inb = 175;
data_ina = 16'h1c0;
data_inb = 16'hffe5;
#10;
address_ina = 176;
address_inb = 177;
data_ina = 16'hfebd;
data_inb = 16'h3ba;
#10;
address_ina = 178;
address_inb = 179;
data_ina = 16'hfc96;
data_inb = 16'hff5e;
#10;
address_ina = 180;
address_inb = 181;
data_ina = 16'hfcad;
data_inb = 16'hfffe;
#10;
address_ina = 182;
address_inb = 183;
data_ina = 16'hfb4c;
data_inb = 16'h644;
#10;
address_ina = 184;
address_inb = 185;
data_ina = 16'hf9d3;
data_inb = 16'hff49;
#10;
address_ina = 186;
address_inb = 187;
data_ina = 16'h3dc;
data_inb = 16'hfae8;
#10;
address_ina = 188;
address_inb = 189;
data_ina = 16'h4d5;
data_inb = 16'hff88;
#10;
address_ina = 190;
address_inb = 191;
data_ina = 16'h37a;
data_inb = 16'h3f2;
#10;
address_ina = 192;
address_inb = 193;
data_ina = 16'h104;
data_inb = 16'h5f1;
#10;
address_ina = 194;
address_inb = 195;
data_ina = 16'hfa87;
data_inb = 16'hff6c;
#10;
address_ina = 196;
address_inb = 197;
data_ina = 16'h429;
data_inb = 16'h1a1;
#10;
address_ina = 198;
address_inb = 199;
data_ina = 16'hffe5;
data_inb = 16'hfcae;
#10;
address_ina = 200;
address_inb = 201;
data_ina = 16'hfd88;
data_inb = 16'h3ad;
#10;
address_ina = 202;
address_inb = 203;
data_ina = 16'hfd13;
data_inb = 16'hff97;
#10;
address_ina = 204;
address_inb = 205;
data_ina = 16'hfec5;
data_inb = 16'hc3;
#10;
address_ina = 206;
address_inb = 207;
data_ina = 16'h42c;
data_inb = 16'hfb68;
#10;
address_ina = 208;
address_inb = 209;
data_ina = 16'h34;
data_inb = 16'h274;
#10;
address_ina = 210;
address_inb = 211;
data_ina = 16'hfca0;
data_inb = 16'h641;
#10;
address_ina = 212;
address_inb = 213;
data_ina = 16'h4c9;
data_inb = 16'h431;
#10;
address_ina = 214;
address_inb = 215;
data_ina = 16'h50b;
data_inb = 16'h669;
#10;
address_ina = 216;
address_inb = 217;
data_ina = 16'hfdaf;
data_inb = 16'h3ec;
#10;
address_ina = 218;
address_inb = 219;
data_ina = 16'h2a3;
data_inb = 16'hfe59;
#10;
address_ina = 220;
address_inb = 221;
data_ina = 16'h332;
data_inb = 16'h11c;
#10;
address_ina = 222;
address_inb = 223;
data_ina = 16'hfa04;
data_inb = 16'h568;
#10;
address_ina = 224;
address_inb = 225;
data_ina = 16'hf9b0;
data_inb = 16'hfd29;
#10;
address_ina = 226;
address_inb = 227;
data_ina = 16'h438;
data_inb = 16'hfee8;
#10;
address_ina = 228;
address_inb = 229;
data_ina = 16'h635;
data_inb = 16'h17d;
#10;
address_ina = 230;
address_inb = 231;
data_ina = 16'hfa0c;
data_inb = 16'h3bc;
#10;
address_ina = 232;
address_inb = 233;
data_ina = 16'hffa7;
data_inb = 16'h49f;
#10;
address_ina = 234;
address_inb = 235;
data_ina = 16'hfacc;
data_inb = 16'hfd00;
#10;
address_ina = 236;
address_inb = 237;
data_ina = 16'h40;
data_inb = 16'hf99c;
#10;
address_ina = 238;
address_inb = 239;
data_ina = 16'hfdec;
data_inb = 16'ha9;
#10;
address_ina = 240;
address_inb = 241;
data_ina = 16'hff07;
data_inb = 16'hffe6;
#10;
address_ina = 242;
address_inb = 243;
data_ina = 16'h613;
data_inb = 16'hfe14;
#10;
address_ina = 244;
address_inb = 245;
data_ina = 16'hfa42;
data_inb = 16'h13d;
#10;
address_ina = 246;
address_inb = 247;
data_ina = 16'h4a;
data_inb = 16'h309;
#10;
address_ina = 248;
address_inb = 249;
data_ina = 16'hf9a4;
data_inb = 16'hfdbb;
#10;
address_ina = 250;
address_inb = 251;
data_ina = 16'hb5;
data_inb = 16'h24c;
#10;
address_ina = 252;
address_inb = 253;
data_ina = 16'h252;
data_inb = 16'h449;
#10;
address_ina = 254;
address_inb = 255;
data_ina = 16'h3d3;
data_inb = 16'hfcc2;
#10;
        wait(init_done);
        #30
        we = 0;
        // Start processing
         
		  #38000

        start = 0;



//        wait (wr_req);
//		  wait (!wr_req);
//		   rd_req = 1;
		  wait(done);
		  #20000
rd_req = 1;
        #70 
		  start = 1;
		 #80 
wait(rd_empty)
rd_req = 0;

$display("Finished the NTT test Number %d",test_num);
////Begin test number #50//////////////
rst = 1;

//#1000
start = 1;
mode = 1; //NTT 0 // INTT 1

// Reset for a few clock cycles

#1000

rst = 0;
test_num = test_num + 1;
#1000
we = 1;
address_ina = 0;
address_inb = 1;
data_ina = 16'hff21;
data_inb = 16'hfa22;
#10;
address_ina = 2;
address_inb = 3;
data_ina = 16'h457;
data_inb = 16'hfecc;
#10;
address_ina = 4;
address_inb = 5;
data_ina = 16'hff3e;
data_inb = 16'hf9ab;
#10;
address_ina = 6;
address_inb = 7;
data_ina = 16'h2c9;
data_inb = 16'hfca2;
#10;
address_ina = 8;
address_inb = 9;
data_ina = 16'hfa45;
data_inb = 16'hfa84;
#10;
address_ina = 10;
address_inb = 11;
data_ina = 16'hfd99;
data_inb = 16'h4ca;
#10;
address_ina = 12;
address_inb = 13;
data_ina = 16'h364;
data_inb = 16'hfb9e;
#10;
address_ina = 14;
address_inb = 15;
data_ina = 16'h4b3;
data_inb = 16'hff77;
#10;
address_ina = 16;
address_inb = 17;
data_ina = 16'h9f;
data_inb = 16'hdc;
#10;
address_ina = 18;
address_inb = 19;
data_ina = 16'hfe5f;
data_inb = 16'hff51;
#10;
address_ina = 20;
address_inb = 21;
data_ina = 16'hfb5e;
data_inb = 16'hfac2;
#10;
address_ina = 22;
address_inb = 23;
data_ina = 16'hff43;
data_inb = 16'h596;
#10;
address_ina = 24;
address_inb = 25;
data_ina = 16'hff94;
data_inb = 16'hfa43;
#10;
address_ina = 26;
address_inb = 27;
data_ina = 16'h14e;
data_inb = 16'hffe2;
#10;
address_ina = 28;
address_inb = 29;
data_ina = 16'hfc8f;
data_inb = 16'h33c;
#10;
address_ina = 30;
address_inb = 31;
data_ina = 16'hfb1f;
data_inb = 16'h12c;
#10;
address_ina = 32;
address_inb = 33;
data_ina = 16'hfdec;
data_inb = 16'hfd50;
#10;
address_ina = 34;
address_inb = 35;
data_ina = 16'hf9b8;
data_inb = 16'h5bc;
#10;
address_ina = 36;
address_inb = 37;
data_ina = 16'hff19;
data_inb = 16'h403;
#10;
address_ina = 38;
address_inb = 39;
data_ina = 16'hfa7f;
data_inb = 16'hff6d;
#10;
address_ina = 40;
address_inb = 41;
data_ina = 16'h53d;
data_inb = 16'hfa1b;
#10;
address_ina = 42;
address_inb = 43;
data_ina = 16'h37;
data_inb = 16'hfa9c;
#10;
address_ina = 44;
address_inb = 45;
data_ina = 16'hfa32;
data_inb = 16'hfe0c;
#10;
address_ina = 46;
address_inb = 47;
data_ina = 16'hfb24;
data_inb = 16'h223;
#10;
address_ina = 48;
address_inb = 49;
data_ina = 16'hfcc0;
data_inb = 16'hffb1;
#10;
address_ina = 50;
address_inb = 51;
data_ina = 16'h48e;
data_inb = 16'h66f;
#10;
address_ina = 52;
address_inb = 53;
data_ina = 16'hfca5;
data_inb = 16'h1a4;
#10;
address_ina = 54;
address_inb = 55;
data_ina = 16'hfd5a;
data_inb = 16'h4d3;
#10;
address_ina = 56;
address_inb = 57;
data_ina = 16'h1d9;
data_inb = 16'h4e6;
#10;
address_ina = 58;
address_inb = 59;
data_ina = 16'hfc6b;
data_inb = 16'hfcb2;
#10;
address_ina = 60;
address_inb = 61;
data_ina = 16'hfdde;
data_inb = 16'hfdd6;
#10;
address_ina = 62;
address_inb = 63;
data_ina = 16'hfcb2;
data_inb = 16'h447;
#10;
address_ina = 64;
address_inb = 65;
data_ina = 16'h350;
data_inb = 16'hfcf4;
#10;
address_ina = 66;
address_inb = 67;
data_ina = 16'hf992;
data_inb = 16'h636;
#10;
address_ina = 68;
address_inb = 69;
data_ina = 16'h32f;
data_inb = 16'hfdb9;
#10;
address_ina = 70;
address_inb = 71;
data_ina = 16'h497;
data_inb = 16'h256;
#10;
address_ina = 72;
address_inb = 73;
data_ina = 16'hfdbe;
data_inb = 16'hfaa5;
#10;
address_ina = 74;
address_inb = 75;
data_ina = 16'hfaa5;
data_inb = 16'hfa40;
#10;
address_ina = 76;
address_inb = 77;
data_ina = 16'h13d;
data_inb = 16'h3e2;
#10;
address_ina = 78;
address_inb = 79;
data_ina = 16'hfdf3;
data_inb = 16'hfc0d;
#10;
address_ina = 80;
address_inb = 81;
data_ina = 16'h5c8;
data_inb = 16'hfc46;
#10;
address_ina = 82;
address_inb = 83;
data_ina = 16'hfa23;
data_inb = 16'h62a;
#10;
address_ina = 84;
address_inb = 85;
data_ina = 16'h3d6;
data_inb = 16'h272;
#10;
address_ina = 86;
address_inb = 87;
data_ina = 16'hfba0;
data_inb = 16'h58b;
#10;
address_ina = 88;
address_inb = 89;
data_ina = 16'hfd23;
data_inb = 16'h63e;
#10;
address_ina = 90;
address_inb = 91;
data_ina = 16'h69;
data_inb = 16'h521;
#10;
address_ina = 92;
address_inb = 93;
data_ina = 16'hbd;
data_inb = 16'hfcdd;
#10;
address_ina = 94;
address_inb = 95;
data_ina = 16'h524;
data_inb = 16'hfb5f;
#10;
address_ina = 96;
address_inb = 97;
data_ina = 16'hfbe0;
data_inb = 16'h5dd;
#10;
address_ina = 98;
address_inb = 99;
data_ina = 16'hfee2;
data_inb = 16'h2f6;
#10;
address_ina = 100;
address_inb = 101;
data_ina = 16'h181;
data_inb = 16'h611;
#10;
address_ina = 102;
address_inb = 103;
data_ina = 16'hff4b;
data_inb = 16'h291;
#10;
address_ina = 104;
address_inb = 105;
data_ina = 16'hf9d9;
data_inb = 16'hfad3;
#10;
address_ina = 106;
address_inb = 107;
data_ina = 16'hfda0;
data_inb = 16'h11;
#10;
address_ina = 108;
address_inb = 109;
data_ina = 16'hff67;
data_inb = 16'hfb80;
#10;
address_ina = 110;
address_inb = 111;
data_ina = 16'h505;
data_inb = 16'h597;
#10;
address_ina = 112;
address_inb = 113;
data_ina = 16'hffe5;
data_inb = 16'hfcb4;
#10;
address_ina = 114;
address_inb = 115;
data_ina = 16'h104;
data_inb = 16'h4c9;
#10;
address_ina = 116;
address_inb = 117;
data_ina = 16'h233;
data_inb = 16'hfccc;
#10;
address_ina = 118;
address_inb = 119;
data_ina = 16'h98;
data_inb = 16'hfab6;
#10;
address_ina = 120;
address_inb = 121;
data_ina = 16'hfe78;
data_inb = 16'h61f;
#10;
address_ina = 122;
address_inb = 123;
data_ina = 16'h182;
data_inb = 16'h1a;
#10;
address_ina = 124;
address_inb = 125;
data_ina = 16'h436;
data_inb = 16'h1b;
#10;
address_ina = 126;
address_inb = 127;
data_ina = 16'h5ce;
data_inb = 16'h498;
#10;
address_ina = 128;
address_inb = 129;
data_ina = 16'h71;
data_inb = 16'hfe4d;
#10;
address_ina = 130;
address_inb = 131;
data_ina = 16'h5a8;
data_inb = 16'h580;
#10;
address_ina = 132;
address_inb = 133;
data_ina = 16'h5bc;
data_inb = 16'h5ca;
#10;
address_ina = 134;
address_inb = 135;
data_ina = 16'hfe17;
data_inb = 16'hfdd0;
#10;
address_ina = 136;
address_inb = 137;
data_ina = 16'h385;
data_inb = 16'hfb32;
#10;
address_ina = 138;
address_inb = 139;
data_ina = 16'hfe63;
data_inb = 16'hf9e8;
#10;
address_ina = 140;
address_inb = 141;
data_ina = 16'h42e;
data_inb = 16'h458;
#10;
address_ina = 142;
address_inb = 143;
data_ina = 16'hff02;
data_inb = 16'hf9a0;
#10;
address_ina = 144;
address_inb = 145;
data_ina = 16'hffb2;
data_inb = 16'hfe18;
#10;
address_ina = 146;
address_inb = 147;
data_ina = 16'hfd9a;
data_inb = 16'h38d;
#10;
address_ina = 148;
address_inb = 149;
data_ina = 16'hfaed;
data_inb = 16'hfb01;
#10;
address_ina = 150;
address_inb = 151;
data_ina = 16'hf9da;
data_inb = 16'h322;
#10;
address_ina = 152;
address_inb = 153;
data_ina = 16'hf9f1;
data_inb = 16'hffd3;
#10;
address_ina = 154;
address_inb = 155;
data_ina = 16'h47c;
data_inb = 16'hfa2b;
#10;
address_ina = 156;
address_inb = 157;
data_ina = 16'h69;
data_inb = 16'h4ee;
#10;
address_ina = 158;
address_inb = 159;
data_ina = 16'hfd7f;
data_inb = 16'hfb14;
#10;
address_ina = 160;
address_inb = 161;
data_ina = 16'hff2e;
data_inb = 16'hfcb6;
#10;
address_ina = 162;
address_inb = 163;
data_ina = 16'hfaf1;
data_inb = 16'hffd8;
#10;
address_ina = 164;
address_inb = 165;
data_ina = 16'hfdeb;
data_inb = 16'hfd29;
#10;
address_ina = 166;
address_inb = 167;
data_ina = 16'h418;
data_inb = 16'ha5;
#10;
address_ina = 168;
address_inb = 169;
data_ina = 16'hfa12;
data_inb = 16'hfbdc;
#10;
address_ina = 170;
address_inb = 171;
data_ina = 16'h4a9;
data_inb = 16'hff9e;
#10;
address_ina = 172;
address_inb = 173;
data_ina = 16'hfdd1;
data_inb = 16'hfa04;
#10;
address_ina = 174;
address_inb = 175;
data_ina = 16'h47a;
data_inb = 16'hff27;
#10;
address_ina = 176;
address_inb = 177;
data_ina = 16'h5f6;
data_inb = 16'h3a;
#10;
address_ina = 178;
address_inb = 179;
data_ina = 16'h20d;
data_inb = 16'hfd8b;
#10;
address_ina = 180;
address_inb = 181;
data_ina = 16'h4c0;
data_inb = 16'hfc7c;
#10;
address_ina = 182;
address_inb = 183;
data_ina = 16'hfd5d;
data_inb = 16'hfa92;
#10;
address_ina = 184;
address_inb = 185;
data_ina = 16'hfb59;
data_inb = 16'hfdf3;
#10;
address_ina = 186;
address_inb = 187;
data_ina = 16'h4f8;
data_inb = 16'hfe9c;
#10;
address_ina = 188;
address_inb = 189;
data_ina = 16'hfbc8;
data_inb = 16'h522;
#10;
address_ina = 190;
address_inb = 191;
data_ina = 16'hfbbc;
data_inb = 16'hff76;
#10;
address_ina = 192;
address_inb = 193;
data_ina = 16'h3d1;
data_inb = 16'h497;
#10;
address_ina = 194;
address_inb = 195;
data_ina = 16'ha3;
data_inb = 16'h17;
#10;
address_ina = 196;
address_inb = 197;
data_ina = 16'h5de;
data_inb = 16'h107;
#10;
address_ina = 198;
address_inb = 199;
data_ina = 16'hfac8;
data_inb = 16'h46c;
#10;
address_ina = 200;
address_inb = 201;
data_ina = 16'hd2;
data_inb = 16'hff1a;
#10;
address_ina = 202;
address_inb = 203;
data_ina = 16'hff0c;
data_inb = 16'hfaa2;
#10;
address_ina = 204;
address_inb = 205;
data_ina = 16'hfef1;
data_inb = 16'he8;
#10;
address_ina = 206;
address_inb = 207;
data_ina = 16'hffba;
data_inb = 16'hc8;
#10;
address_ina = 208;
address_inb = 209;
data_ina = 16'hfedd;
data_inb = 16'h158;
#10;
address_ina = 210;
address_inb = 211;
data_ina = 16'h63c;
data_inb = 16'hd6;
#10;
address_ina = 212;
address_inb = 213;
data_ina = 16'h4ae;
data_inb = 16'hfd17;
#10;
address_ina = 214;
address_inb = 215;
data_ina = 16'h137;
data_inb = 16'hf9b4;
#10;
address_ina = 216;
address_inb = 217;
data_ina = 16'hfda5;
data_inb = 16'hf99c;
#10;
address_ina = 218;
address_inb = 219;
data_ina = 16'h7c;
data_inb = 16'h62f;
#10;
address_ina = 220;
address_inb = 221;
data_ina = 16'h1e3;
data_inb = 16'hf99a;
#10;
address_ina = 222;
address_inb = 223;
data_ina = 16'h178;
data_inb = 16'hfd83;
#10;
address_ina = 224;
address_inb = 225;
data_ina = 16'he9;
data_inb = 16'h627;
#10;
address_ina = 226;
address_inb = 227;
data_ina = 16'hf9db;
data_inb = 16'ha8;
#10;
address_ina = 228;
address_inb = 229;
data_ina = 16'hfd0e;
data_inb = 16'h24a;
#10;
address_ina = 230;
address_inb = 231;
data_ina = 16'hfe5c;
data_inb = 16'h2e2;
#10;
address_ina = 232;
address_inb = 233;
data_ina = 16'hfb28;
data_inb = 16'h55f;
#10;
address_ina = 234;
address_inb = 235;
data_ina = 16'h23b;
data_inb = 16'hf980;
#10;
address_ina = 236;
address_inb = 237;
data_ina = 16'hfb33;
data_inb = 16'hfe36;
#10;
address_ina = 238;
address_inb = 239;
data_ina = 16'h154;
data_inb = 16'h66b;
#10;
address_ina = 240;
address_inb = 241;
data_ina = 16'hff78;
data_inb = 16'h2f;
#10;
address_ina = 242;
address_inb = 243;
data_ina = 16'h60a;
data_inb = 16'hfd43;
#10;
address_ina = 244;
address_inb = 245;
data_ina = 16'h7c;
data_inb = 16'h4ed;
#10;
address_ina = 246;
address_inb = 247;
data_ina = 16'hff7c;
data_inb = 16'h74;
#10;
address_ina = 248;
address_inb = 249;
data_ina = 16'h1fd;
data_inb = 16'hfab9;
#10;
address_ina = 250;
address_inb = 251;
data_ina = 16'hfb9a;
data_inb = 16'hff50;
#10;
address_ina = 252;
address_inb = 253;
data_ina = 16'h610;
data_inb = 16'hfa1a;
#10;
address_ina = 254;
address_inb = 255;
data_ina = 16'hff0c;
data_inb = 16'h494;
#10;
        wait(init_done);
        #30
        we = 0;
        // Start processing
         
		  #38000

        start = 0;



//        wait (wr_req);
//		  wait (!wr_req);
//		   rd_req = 1;
		  wait(done);
		  #20000
rd_req = 1;
        #70 
		  start = 1;
		 #80 
wait(rd_empty)
rd_req = 0;

$display("Finished the NTT test Number %d",test_num);
////Begin test number #51//////////////
rst = 1;

//#1000
start = 1;
mode = 0; //NTT 0 // INTT 1

// Reset for a few clock cycles

#1000

rst = 0;
test_num = test_num + 1;
#1000
we = 1;
address_ina = 0;
address_inb = 1;
data_ina = 16'hfffe;
data_inb = 16'h0;
#10;
address_ina = 2;
address_inb = 3;
data_ina = 16'h0;
data_inb = 16'hfffe;
#10;
address_ina = 4;
address_inb = 5;
data_ina = 16'h3;
data_inb = 16'h0;
#10;
address_ina = 6;
address_inb = 7;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 8;
address_inb = 9;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 10;
address_inb = 11;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 12;
address_inb = 13;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 14;
address_inb = 15;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 16;
address_inb = 17;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 18;
address_inb = 19;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 20;
address_inb = 21;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 22;
address_inb = 23;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 24;
address_inb = 25;
data_ina = 16'h1;
data_inb = 16'hfffd;
#10;
address_ina = 26;
address_inb = 27;
data_ina = 16'h2;
data_inb = 16'hfffe;
#10;
address_ina = 28;
address_inb = 29;
data_ina = 16'h0;
data_inb = 16'hfffe;
#10;
address_ina = 30;
address_inb = 31;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 32;
address_inb = 33;
data_ina = 16'hfffe;
data_inb = 16'h0;
#10;
address_ina = 34;
address_inb = 35;
data_ina = 16'h2;
data_inb = 16'h3;
#10;
address_ina = 36;
address_inb = 37;
data_ina = 16'h3;
data_inb = 16'h0;
#10;
address_ina = 38;
address_inb = 39;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 40;
address_inb = 41;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 42;
address_inb = 43;
data_ina = 16'h2;
data_inb = 16'hfffe;
#10;
address_ina = 44;
address_inb = 45;
data_ina = 16'h2;
data_inb = 16'hffff;
#10;
address_ina = 46;
address_inb = 47;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 48;
address_inb = 49;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 50;
address_inb = 51;
data_ina = 16'hfffe;
data_inb = 16'h0;
#10;
address_ina = 52;
address_inb = 53;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 54;
address_inb = 55;
data_ina = 16'h0;
data_inb = 16'h3;
#10;
address_ina = 56;
address_inb = 57;
data_ina = 16'hfffe;
data_inb = 16'hffff;
#10;
address_ina = 58;
address_inb = 59;
data_ina = 16'h1;
data_inb = 16'h2;
#10;
address_ina = 60;
address_inb = 61;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 62;
address_inb = 63;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 64;
address_inb = 65;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 66;
address_inb = 67;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 68;
address_inb = 69;
data_ina = 16'h2;
data_inb = 16'hffff;
#10;
address_ina = 70;
address_inb = 71;
data_ina = 16'h0;
data_inb = 16'hfffe;
#10;
address_ina = 72;
address_inb = 73;
data_ina = 16'hfffe;
data_inb = 16'hffff;
#10;
address_ina = 74;
address_inb = 75;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 76;
address_inb = 77;
data_ina = 16'hfffe;
data_inb = 16'h0;
#10;
address_ina = 78;
address_inb = 79;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 80;
address_inb = 81;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 82;
address_inb = 83;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 84;
address_inb = 85;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 86;
address_inb = 87;
data_ina = 16'h2;
data_inb = 16'h1;
#10;
address_ina = 88;
address_inb = 89;
data_ina = 16'h1;
data_inb = 16'hfffe;
#10;
address_ina = 90;
address_inb = 91;
data_ina = 16'h2;
data_inb = 16'h2;
#10;
address_ina = 92;
address_inb = 93;
data_ina = 16'h1;
data_inb = 16'hfffe;
#10;
address_ina = 94;
address_inb = 95;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 96;
address_inb = 97;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 98;
address_inb = 99;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 100;
address_inb = 101;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 102;
address_inb = 103;
data_ina = 16'hffff;
data_inb = 16'hfffe;
#10;
address_ina = 104;
address_inb = 105;
data_ina = 16'hfffd;
data_inb = 16'hfffe;
#10;
address_ina = 106;
address_inb = 107;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 108;
address_inb = 109;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 110;
address_inb = 111;
data_ina = 16'hfffd;
data_inb = 16'h0;
#10;
address_ina = 112;
address_inb = 113;
data_ina = 16'h2;
data_inb = 16'hfffe;
#10;
address_ina = 114;
address_inb = 115;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 116;
address_inb = 117;
data_ina = 16'hfffe;
data_inb = 16'h0;
#10;
address_ina = 118;
address_inb = 119;
data_ina = 16'hfffe;
data_inb = 16'h0;
#10;
address_ina = 120;
address_inb = 121;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 122;
address_inb = 123;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 124;
address_inb = 125;
data_ina = 16'hfffe;
data_inb = 16'h1;
#10;
address_ina = 126;
address_inb = 127;
data_ina = 16'hfffe;
data_inb = 16'h0;
#10;
address_ina = 128;
address_inb = 129;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 130;
address_inb = 131;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 132;
address_inb = 133;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 134;
address_inb = 135;
data_ina = 16'h2;
data_inb = 16'h1;
#10;
address_ina = 136;
address_inb = 137;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 138;
address_inb = 139;
data_ina = 16'h2;
data_inb = 16'h2;
#10;
address_ina = 140;
address_inb = 141;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 142;
address_inb = 143;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 144;
address_inb = 145;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 146;
address_inb = 147;
data_ina = 16'h2;
data_inb = 16'hffff;
#10;
address_ina = 148;
address_inb = 149;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 150;
address_inb = 151;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 152;
address_inb = 153;
data_ina = 16'h2;
data_inb = 16'hfffe;
#10;
address_ina = 154;
address_inb = 155;
data_ina = 16'h1;
data_inb = 16'h2;
#10;
address_ina = 156;
address_inb = 157;
data_ina = 16'hffff;
data_inb = 16'hfffe;
#10;
address_ina = 158;
address_inb = 159;
data_ina = 16'hffff;
data_inb = 16'hfffe;
#10;
address_ina = 160;
address_inb = 161;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 162;
address_inb = 163;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 164;
address_inb = 165;
data_ina = 16'hffff;
data_inb = 16'hfffe;
#10;
address_ina = 166;
address_inb = 167;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 168;
address_inb = 169;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 170;
address_inb = 171;
data_ina = 16'hfffe;
data_inb = 16'hffff;
#10;
address_ina = 172;
address_inb = 173;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 174;
address_inb = 175;
data_ina = 16'h2;
data_inb = 16'hffff;
#10;
address_ina = 176;
address_inb = 177;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 178;
address_inb = 179;
data_ina = 16'hfffe;
data_inb = 16'h0;
#10;
address_ina = 180;
address_inb = 181;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 182;
address_inb = 183;
data_ina = 16'h1;
data_inb = 16'h2;
#10;
address_ina = 184;
address_inb = 185;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 186;
address_inb = 187;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 188;
address_inb = 189;
data_ina = 16'h0;
data_inb = 16'hfffe;
#10;
address_ina = 190;
address_inb = 191;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 192;
address_inb = 193;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 194;
address_inb = 195;
data_ina = 16'h0;
data_inb = 16'h2;
#10;
address_ina = 196;
address_inb = 197;
data_ina = 16'h0;
data_inb = 16'h2;
#10;
address_ina = 198;
address_inb = 199;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 200;
address_inb = 201;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 202;
address_inb = 203;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 204;
address_inb = 205;
data_ina = 16'hfffe;
data_inb = 16'hfffe;
#10;
address_ina = 206;
address_inb = 207;
data_ina = 16'hffff;
data_inb = 16'hfffe;
#10;
address_ina = 208;
address_inb = 209;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 210;
address_inb = 211;
data_ina = 16'hfffe;
data_inb = 16'h0;
#10;
address_ina = 212;
address_inb = 213;
data_ina = 16'hfffe;
data_inb = 16'hffff;
#10;
address_ina = 214;
address_inb = 215;
data_ina = 16'hfffd;
data_inb = 16'hfffe;
#10;
address_ina = 216;
address_inb = 217;
data_ina = 16'h1;
data_inb = 16'hfffe;
#10;
address_ina = 218;
address_inb = 219;
data_ina = 16'hfffe;
data_inb = 16'h0;
#10;
address_ina = 220;
address_inb = 221;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 222;
address_inb = 223;
data_ina = 16'h0;
data_inb = 16'h2;
#10;
address_ina = 224;
address_inb = 225;
data_ina = 16'hfffe;
data_inb = 16'h2;
#10;
address_ina = 226;
address_inb = 227;
data_ina = 16'h0;
data_inb = 16'hfffe;
#10;
address_ina = 228;
address_inb = 229;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 230;
address_inb = 231;
data_ina = 16'hffff;
data_inb = 16'hfffe;
#10;
address_ina = 232;
address_inb = 233;
data_ina = 16'hfffe;
data_inb = 16'hffff;
#10;
address_ina = 234;
address_inb = 235;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 236;
address_inb = 237;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 238;
address_inb = 239;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 240;
address_inb = 241;
data_ina = 16'h0;
data_inb = 16'h2;
#10;
address_ina = 242;
address_inb = 243;
data_ina = 16'hfffe;
data_inb = 16'h1;
#10;
address_ina = 244;
address_inb = 245;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 246;
address_inb = 247;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 248;
address_inb = 249;
data_ina = 16'h1;
data_inb = 16'hfffe;
#10;
address_ina = 250;
address_inb = 251;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 252;
address_inb = 253;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 254;
address_inb = 255;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
        wait(init_done);
        #30
        we = 0;
        // Start processing
         
		  #38000

        start = 0;



//        wait (wr_req);
//		  wait (!wr_req);
//		   rd_req = 1;
		  wait(done);
		  #20000
rd_req = 1;
        #70 
		  start = 1;
		 #80 
wait(rd_empty)
rd_req = 0;

$display("Finished the NTT test Number %d",test_num);
////Begin test number #52//////////////
rst = 1;

//#1000
start = 1;
mode = 0; //NTT 0 // INTT 1

// Reset for a few clock cycles

#1000

rst = 0;
test_num = test_num + 1;
#1000
we = 1;
address_ina = 0;
address_inb = 1;
data_ina = 16'h2;
data_inb = 16'hffff;
#10;
address_ina = 2;
address_inb = 3;
data_ina = 16'hfffd;
data_inb = 16'h0;
#10;
address_ina = 4;
address_inb = 5;
data_ina = 16'h2;
data_inb = 16'hfffe;
#10;
address_ina = 6;
address_inb = 7;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 8;
address_inb = 9;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 10;
address_inb = 11;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 12;
address_inb = 13;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 14;
address_inb = 15;
data_ina = 16'hfffe;
data_inb = 16'h1;
#10;
address_ina = 16;
address_inb = 17;
data_ina = 16'h1;
data_inb = 16'hfffe;
#10;
address_ina = 18;
address_inb = 19;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 20;
address_inb = 21;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 22;
address_inb = 23;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 24;
address_inb = 25;
data_ina = 16'hfffe;
data_inb = 16'hffff;
#10;
address_ina = 26;
address_inb = 27;
data_ina = 16'h0;
data_inb = 16'hfffe;
#10;
address_ina = 28;
address_inb = 29;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 30;
address_inb = 31;
data_ina = 16'h1;
data_inb = 16'hfffe;
#10;
address_ina = 32;
address_inb = 33;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 34;
address_inb = 35;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 36;
address_inb = 37;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 38;
address_inb = 39;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 40;
address_inb = 41;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 42;
address_inb = 43;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 44;
address_inb = 45;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 46;
address_inb = 47;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 48;
address_inb = 49;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 50;
address_inb = 51;
data_ina = 16'h0;
data_inb = 16'hfffe;
#10;
address_ina = 52;
address_inb = 53;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 54;
address_inb = 55;
data_ina = 16'hfffe;
data_inb = 16'hfffe;
#10;
address_ina = 56;
address_inb = 57;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 58;
address_inb = 59;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 60;
address_inb = 61;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 62;
address_inb = 63;
data_ina = 16'h2;
data_inb = 16'h1;
#10;
address_ina = 64;
address_inb = 65;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 66;
address_inb = 67;
data_ina = 16'h0;
data_inb = 16'hfffe;
#10;
address_ina = 68;
address_inb = 69;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 70;
address_inb = 71;
data_ina = 16'hfffe;
data_inb = 16'hfffe;
#10;
address_ina = 72;
address_inb = 73;
data_ina = 16'hfffe;
data_inb = 16'hffff;
#10;
address_ina = 74;
address_inb = 75;
data_ina = 16'h2;
data_inb = 16'h1;
#10;
address_ina = 76;
address_inb = 77;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 78;
address_inb = 79;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 80;
address_inb = 81;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 82;
address_inb = 83;
data_ina = 16'h2;
data_inb = 16'h0;
#10;
address_ina = 84;
address_inb = 85;
data_ina = 16'hfffe;
data_inb = 16'hffff;
#10;
address_ina = 86;
address_inb = 87;
data_ina = 16'hfffe;
data_inb = 16'hffff;
#10;
address_ina = 88;
address_inb = 89;
data_ina = 16'hfffe;
data_inb = 16'hffff;
#10;
address_ina = 90;
address_inb = 91;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 92;
address_inb = 93;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 94;
address_inb = 95;
data_ina = 16'h2;
data_inb = 16'h2;
#10;
address_ina = 96;
address_inb = 97;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 98;
address_inb = 99;
data_ina = 16'hfffd;
data_inb = 16'h0;
#10;
address_ina = 100;
address_inb = 101;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 102;
address_inb = 103;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 104;
address_inb = 105;
data_ina = 16'h1;
data_inb = 16'h3;
#10;
address_ina = 106;
address_inb = 107;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 108;
address_inb = 109;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 110;
address_inb = 111;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 112;
address_inb = 113;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 114;
address_inb = 115;
data_ina = 16'h1;
data_inb = 16'hfffe;
#10;
address_ina = 116;
address_inb = 117;
data_ina = 16'h0;
data_inb = 16'h2;
#10;
address_ina = 118;
address_inb = 119;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 120;
address_inb = 121;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 122;
address_inb = 123;
data_ina = 16'h0;
data_inb = 16'h3;
#10;
address_ina = 124;
address_inb = 125;
data_ina = 16'h2;
data_inb = 16'h2;
#10;
address_ina = 126;
address_inb = 127;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 128;
address_inb = 129;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 130;
address_inb = 131;
data_ina = 16'h1;
data_inb = 16'h2;
#10;
address_ina = 132;
address_inb = 133;
data_ina = 16'h0;
data_inb = 16'h2;
#10;
address_ina = 134;
address_inb = 135;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 136;
address_inb = 137;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 138;
address_inb = 139;
data_ina = 16'h2;
data_inb = 16'h0;
#10;
address_ina = 140;
address_inb = 141;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 142;
address_inb = 143;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 144;
address_inb = 145;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 146;
address_inb = 147;
data_ina = 16'hffff;
data_inb = 16'h3;
#10;
address_ina = 148;
address_inb = 149;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 150;
address_inb = 151;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 152;
address_inb = 153;
data_ina = 16'h1;
data_inb = 16'h2;
#10;
address_ina = 154;
address_inb = 155;
data_ina = 16'hfffe;
data_inb = 16'h0;
#10;
address_ina = 156;
address_inb = 157;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 158;
address_inb = 159;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 160;
address_inb = 161;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 162;
address_inb = 163;
data_ina = 16'hfffe;
data_inb = 16'h1;
#10;
address_ina = 164;
address_inb = 165;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 166;
address_inb = 167;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 168;
address_inb = 169;
data_ina = 16'h1;
data_inb = 16'hfffe;
#10;
address_ina = 170;
address_inb = 171;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 172;
address_inb = 173;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 174;
address_inb = 175;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 176;
address_inb = 177;
data_ina = 16'hfffe;
data_inb = 16'h0;
#10;
address_ina = 178;
address_inb = 179;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 180;
address_inb = 181;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 182;
address_inb = 183;
data_ina = 16'h2;
data_inb = 16'h0;
#10;
address_ina = 184;
address_inb = 185;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 186;
address_inb = 187;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 188;
address_inb = 189;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 190;
address_inb = 191;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 192;
address_inb = 193;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 194;
address_inb = 195;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 196;
address_inb = 197;
data_ina = 16'h2;
data_inb = 16'hfffd;
#10;
address_ina = 198;
address_inb = 199;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 200;
address_inb = 201;
data_ina = 16'h1;
data_inb = 16'h2;
#10;
address_ina = 202;
address_inb = 203;
data_ina = 16'hfffe;
data_inb = 16'h0;
#10;
address_ina = 204;
address_inb = 205;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 206;
address_inb = 207;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 208;
address_inb = 209;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 210;
address_inb = 211;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 212;
address_inb = 213;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 214;
address_inb = 215;
data_ina = 16'hfffe;
data_inb = 16'h1;
#10;
address_ina = 216;
address_inb = 217;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 218;
address_inb = 219;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 220;
address_inb = 221;
data_ina = 16'h1;
data_inb = 16'h2;
#10;
address_ina = 222;
address_inb = 223;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 224;
address_inb = 225;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 226;
address_inb = 227;
data_ina = 16'hffff;
data_inb = 16'h2;
#10;
address_ina = 228;
address_inb = 229;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 230;
address_inb = 231;
data_ina = 16'hfffe;
data_inb = 16'h0;
#10;
address_ina = 232;
address_inb = 233;
data_ina = 16'hffff;
data_inb = 16'h2;
#10;
address_ina = 234;
address_inb = 235;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 236;
address_inb = 237;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 238;
address_inb = 239;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 240;
address_inb = 241;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 242;
address_inb = 243;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 244;
address_inb = 245;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 246;
address_inb = 247;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 248;
address_inb = 249;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 250;
address_inb = 251;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 252;
address_inb = 253;
data_ina = 16'hffff;
data_inb = 16'h2;
#10;
address_ina = 254;
address_inb = 255;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
        wait(init_done);
        #30
        we = 0;
        // Start processing
         
		  #38000

        start = 0;



//        wait (wr_req);
//		  wait (!wr_req);
//		   rd_req = 1;
		  wait(done);
		  #20000
rd_req = 1;
        #70 
		  start = 1;
		 #80 
wait(rd_empty)
rd_req = 0;

$display("Finished the NTT test Number %d",test_num);
////Begin test number #53//////////////
rst = 1;

//#1000
start = 1;
mode = 0; //NTT 0 // INTT 1

// Reset for a few clock cycles

#1000

rst = 0;
test_num = test_num + 1;
#1000
we = 1;
address_ina = 0;
address_inb = 1;
data_ina = 16'h2;
data_inb = 16'h0;
#10;
address_ina = 2;
address_inb = 3;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 4;
address_inb = 5;
data_ina = 16'h2;
data_inb = 16'h2;
#10;
address_ina = 6;
address_inb = 7;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 8;
address_inb = 9;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 10;
address_inb = 11;
data_ina = 16'h0;
data_inb = 16'h2;
#10;
address_ina = 12;
address_inb = 13;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 14;
address_inb = 15;
data_ina = 16'hfffe;
data_inb = 16'h1;
#10;
address_ina = 16;
address_inb = 17;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 18;
address_inb = 19;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 20;
address_inb = 21;
data_ina = 16'hfffe;
data_inb = 16'h1;
#10;
address_ina = 22;
address_inb = 23;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 24;
address_inb = 25;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 26;
address_inb = 27;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 28;
address_inb = 29;
data_ina = 16'hffff;
data_inb = 16'h2;
#10;
address_ina = 30;
address_inb = 31;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 32;
address_inb = 33;
data_ina = 16'h2;
data_inb = 16'h0;
#10;
address_ina = 34;
address_inb = 35;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 36;
address_inb = 37;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 38;
address_inb = 39;
data_ina = 16'hfffe;
data_inb = 16'h1;
#10;
address_ina = 40;
address_inb = 41;
data_ina = 16'h1;
data_inb = 16'hfffd;
#10;
address_ina = 42;
address_inb = 43;
data_ina = 16'hfffe;
data_inb = 16'h0;
#10;
address_ina = 44;
address_inb = 45;
data_ina = 16'h0;
data_inb = 16'h2;
#10;
address_ina = 46;
address_inb = 47;
data_ina = 16'hfffe;
data_inb = 16'h0;
#10;
address_ina = 48;
address_inb = 49;
data_ina = 16'h0;
data_inb = 16'hfffe;
#10;
address_ina = 50;
address_inb = 51;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 52;
address_inb = 53;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 54;
address_inb = 55;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 56;
address_inb = 57;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 58;
address_inb = 59;
data_ina = 16'hfffe;
data_inb = 16'h0;
#10;
address_ina = 60;
address_inb = 61;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 62;
address_inb = 63;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 64;
address_inb = 65;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 66;
address_inb = 67;
data_ina = 16'hfffe;
data_inb = 16'h0;
#10;
address_ina = 68;
address_inb = 69;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 70;
address_inb = 71;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 72;
address_inb = 73;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 74;
address_inb = 75;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 76;
address_inb = 77;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 78;
address_inb = 79;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 80;
address_inb = 81;
data_ina = 16'h2;
data_inb = 16'hffff;
#10;
address_ina = 82;
address_inb = 83;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 84;
address_inb = 85;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 86;
address_inb = 87;
data_ina = 16'hfffe;
data_inb = 16'hffff;
#10;
address_ina = 88;
address_inb = 89;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 90;
address_inb = 91;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 92;
address_inb = 93;
data_ina = 16'hffff;
data_inb = 16'h2;
#10;
address_ina = 94;
address_inb = 95;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 96;
address_inb = 97;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 98;
address_inb = 99;
data_ina = 16'h3;
data_inb = 16'hffff;
#10;
address_ina = 100;
address_inb = 101;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 102;
address_inb = 103;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 104;
address_inb = 105;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 106;
address_inb = 107;
data_ina = 16'hfffe;
data_inb = 16'hffff;
#10;
address_ina = 108;
address_inb = 109;
data_ina = 16'h0;
data_inb = 16'hfffe;
#10;
address_ina = 110;
address_inb = 111;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 112;
address_inb = 113;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 114;
address_inb = 115;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 116;
address_inb = 117;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 118;
address_inb = 119;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 120;
address_inb = 121;
data_ina = 16'h1;
data_inb = 16'hfffe;
#10;
address_ina = 122;
address_inb = 123;
data_ina = 16'h2;
data_inb = 16'h0;
#10;
address_ina = 124;
address_inb = 125;
data_ina = 16'h2;
data_inb = 16'hfffe;
#10;
address_ina = 126;
address_inb = 127;
data_ina = 16'hfffe;
data_inb = 16'hfffe;
#10;
address_ina = 128;
address_inb = 129;
data_ina = 16'h2;
data_inb = 16'hffff;
#10;
address_ina = 130;
address_inb = 131;
data_ina = 16'hffff;
data_inb = 16'h3;
#10;
address_ina = 132;
address_inb = 133;
data_ina = 16'h3;
data_inb = 16'h2;
#10;
address_ina = 134;
address_inb = 135;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 136;
address_inb = 137;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 138;
address_inb = 139;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 140;
address_inb = 141;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 142;
address_inb = 143;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 144;
address_inb = 145;
data_ina = 16'h0;
data_inb = 16'hfffe;
#10;
address_ina = 146;
address_inb = 147;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 148;
address_inb = 149;
data_ina = 16'h0;
data_inb = 16'h2;
#10;
address_ina = 150;
address_inb = 151;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 152;
address_inb = 153;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 154;
address_inb = 155;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 156;
address_inb = 157;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 158;
address_inb = 159;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 160;
address_inb = 161;
data_ina = 16'hffff;
data_inb = 16'hfffe;
#10;
address_ina = 162;
address_inb = 163;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 164;
address_inb = 165;
data_ina = 16'h0;
data_inb = 16'hfffe;
#10;
address_ina = 166;
address_inb = 167;
data_ina = 16'hfffe;
data_inb = 16'h0;
#10;
address_ina = 168;
address_inb = 169;
data_ina = 16'h0;
data_inb = 16'h2;
#10;
address_ina = 170;
address_inb = 171;
data_ina = 16'h2;
data_inb = 16'h0;
#10;
address_ina = 172;
address_inb = 173;
data_ina = 16'h1;
data_inb = 16'hfffe;
#10;
address_ina = 174;
address_inb = 175;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 176;
address_inb = 177;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 178;
address_inb = 179;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 180;
address_inb = 181;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 182;
address_inb = 183;
data_ina = 16'h0;
data_inb = 16'h2;
#10;
address_ina = 184;
address_inb = 185;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 186;
address_inb = 187;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 188;
address_inb = 189;
data_ina = 16'hfffe;
data_inb = 16'hfffd;
#10;
address_ina = 190;
address_inb = 191;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 192;
address_inb = 193;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 194;
address_inb = 195;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 196;
address_inb = 197;
data_ina = 16'h1;
data_inb = 16'hfffe;
#10;
address_ina = 198;
address_inb = 199;
data_ina = 16'hfffd;
data_inb = 16'h1;
#10;
address_ina = 200;
address_inb = 201;
data_ina = 16'hfffd;
data_inb = 16'h0;
#10;
address_ina = 202;
address_inb = 203;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 204;
address_inb = 205;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 206;
address_inb = 207;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 208;
address_inb = 209;
data_ina = 16'h2;
data_inb = 16'hffff;
#10;
address_ina = 210;
address_inb = 211;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 212;
address_inb = 213;
data_ina = 16'hfffe;
data_inb = 16'h1;
#10;
address_ina = 214;
address_inb = 215;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 216;
address_inb = 217;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 218;
address_inb = 219;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 220;
address_inb = 221;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 222;
address_inb = 223;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 224;
address_inb = 225;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 226;
address_inb = 227;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 228;
address_inb = 229;
data_ina = 16'hfffe;
data_inb = 16'h0;
#10;
address_ina = 230;
address_inb = 231;
data_ina = 16'hfffe;
data_inb = 16'hffff;
#10;
address_ina = 232;
address_inb = 233;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 234;
address_inb = 235;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 236;
address_inb = 237;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 238;
address_inb = 239;
data_ina = 16'h0;
data_inb = 16'hfffe;
#10;
address_ina = 240;
address_inb = 241;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 242;
address_inb = 243;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 244;
address_inb = 245;
data_ina = 16'h0;
data_inb = 16'h2;
#10;
address_ina = 246;
address_inb = 247;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 248;
address_inb = 249;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 250;
address_inb = 251;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 252;
address_inb = 253;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 254;
address_inb = 255;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
        wait(init_done);
        #30
        we = 0;
        // Start processing
         
		  #38000

        start = 0;



//        wait (wr_req);
//		  wait (!wr_req);
//		   rd_req = 1;
		  wait(done);
		  #20000
rd_req = 1;
        #70 
		  start = 1;
		 #80 
wait(rd_empty)
rd_req = 0;

$display("Finished the NTT test Number %d",test_num);
////Begin test number #54//////////////
rst = 1;

//#1000
start = 1;
mode = 0; //NTT 0 // INTT 1

// Reset for a few clock cycles

#1000

rst = 0;
test_num = test_num + 1;
#1000
we = 1;
address_ina = 0;
address_inb = 1;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 2;
address_inb = 3;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 4;
address_inb = 5;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 6;
address_inb = 7;
data_ina = 16'h1;
data_inb = 16'h2;
#10;
address_ina = 8;
address_inb = 9;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 10;
address_inb = 11;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 12;
address_inb = 13;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 14;
address_inb = 15;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 16;
address_inb = 17;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 18;
address_inb = 19;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 20;
address_inb = 21;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 22;
address_inb = 23;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 24;
address_inb = 25;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 26;
address_inb = 27;
data_ina = 16'h2;
data_inb = 16'hffff;
#10;
address_ina = 28;
address_inb = 29;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 30;
address_inb = 31;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 32;
address_inb = 33;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 34;
address_inb = 35;
data_ina = 16'h2;
data_inb = 16'h1;
#10;
address_ina = 36;
address_inb = 37;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 38;
address_inb = 39;
data_ina = 16'hfffe;
data_inb = 16'h2;
#10;
address_ina = 40;
address_inb = 41;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 42;
address_inb = 43;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 44;
address_inb = 45;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 46;
address_inb = 47;
data_ina = 16'hfffe;
data_inb = 16'h1;
#10;
address_ina = 48;
address_inb = 49;
data_ina = 16'hfffe;
data_inb = 16'h1;
#10;
address_ina = 50;
address_inb = 51;
data_ina = 16'h0;
data_inb = 16'hfffe;
#10;
address_ina = 52;
address_inb = 53;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 54;
address_inb = 55;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 56;
address_inb = 57;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 58;
address_inb = 59;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 60;
address_inb = 61;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 62;
address_inb = 63;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 64;
address_inb = 65;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 66;
address_inb = 67;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 68;
address_inb = 69;
data_ina = 16'h0;
data_inb = 16'hfffe;
#10;
address_ina = 70;
address_inb = 71;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 72;
address_inb = 73;
data_ina = 16'hfffe;
data_inb = 16'h2;
#10;
address_ina = 74;
address_inb = 75;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 76;
address_inb = 77;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 78;
address_inb = 79;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 80;
address_inb = 81;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 82;
address_inb = 83;
data_ina = 16'hffff;
data_inb = 16'hfffe;
#10;
address_ina = 84;
address_inb = 85;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 86;
address_inb = 87;
data_ina = 16'h1;
data_inb = 16'hfffe;
#10;
address_ina = 88;
address_inb = 89;
data_ina = 16'h3;
data_inb = 16'h1;
#10;
address_ina = 90;
address_inb = 91;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 92;
address_inb = 93;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 94;
address_inb = 95;
data_ina = 16'h0;
data_inb = 16'h2;
#10;
address_ina = 96;
address_inb = 97;
data_ina = 16'hfffe;
data_inb = 16'h2;
#10;
address_ina = 98;
address_inb = 99;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 100;
address_inb = 101;
data_ina = 16'h1;
data_inb = 16'hfffd;
#10;
address_ina = 102;
address_inb = 103;
data_ina = 16'h1;
data_inb = 16'h2;
#10;
address_ina = 104;
address_inb = 105;
data_ina = 16'h2;
data_inb = 16'h1;
#10;
address_ina = 106;
address_inb = 107;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 108;
address_inb = 109;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 110;
address_inb = 111;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 112;
address_inb = 113;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 114;
address_inb = 115;
data_ina = 16'h3;
data_inb = 16'h0;
#10;
address_ina = 116;
address_inb = 117;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 118;
address_inb = 119;
data_ina = 16'hffff;
data_inb = 16'h2;
#10;
address_ina = 120;
address_inb = 121;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 122;
address_inb = 123;
data_ina = 16'hfffe;
data_inb = 16'hffff;
#10;
address_ina = 124;
address_inb = 125;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 126;
address_inb = 127;
data_ina = 16'h3;
data_inb = 16'h3;
#10;
address_ina = 128;
address_inb = 129;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 130;
address_inb = 131;
data_ina = 16'hfffe;
data_inb = 16'h2;
#10;
address_ina = 132;
address_inb = 133;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 134;
address_inb = 135;
data_ina = 16'h1;
data_inb = 16'h2;
#10;
address_ina = 136;
address_inb = 137;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 138;
address_inb = 139;
data_ina = 16'h2;
data_inb = 16'hffff;
#10;
address_ina = 140;
address_inb = 141;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 142;
address_inb = 143;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 144;
address_inb = 145;
data_ina = 16'h2;
data_inb = 16'h2;
#10;
address_ina = 146;
address_inb = 147;
data_ina = 16'hfffe;
data_inb = 16'h1;
#10;
address_ina = 148;
address_inb = 149;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 150;
address_inb = 151;
data_ina = 16'hffff;
data_inb = 16'h2;
#10;
address_ina = 152;
address_inb = 153;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 154;
address_inb = 155;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 156;
address_inb = 157;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 158;
address_inb = 159;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 160;
address_inb = 161;
data_ina = 16'hfffe;
data_inb = 16'hffff;
#10;
address_ina = 162;
address_inb = 163;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 164;
address_inb = 165;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 166;
address_inb = 167;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 168;
address_inb = 169;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 170;
address_inb = 171;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 172;
address_inb = 173;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 174;
address_inb = 175;
data_ina = 16'h0;
data_inb = 16'h2;
#10;
address_ina = 176;
address_inb = 177;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 178;
address_inb = 179;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 180;
address_inb = 181;
data_ina = 16'h0;
data_inb = 16'hfffe;
#10;
address_ina = 182;
address_inb = 183;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 184;
address_inb = 185;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 186;
address_inb = 187;
data_ina = 16'hffff;
data_inb = 16'h2;
#10;
address_ina = 188;
address_inb = 189;
data_ina = 16'hfffe;
data_inb = 16'h1;
#10;
address_ina = 190;
address_inb = 191;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 192;
address_inb = 193;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 194;
address_inb = 195;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 196;
address_inb = 197;
data_ina = 16'h3;
data_inb = 16'hfffe;
#10;
address_ina = 198;
address_inb = 199;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 200;
address_inb = 201;
data_ina = 16'h1;
data_inb = 16'h2;
#10;
address_ina = 202;
address_inb = 203;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 204;
address_inb = 205;
data_ina = 16'h0;
data_inb = 16'h2;
#10;
address_ina = 206;
address_inb = 207;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 208;
address_inb = 209;
data_ina = 16'h3;
data_inb = 16'h2;
#10;
address_ina = 210;
address_inb = 211;
data_ina = 16'h1;
data_inb = 16'h2;
#10;
address_ina = 212;
address_inb = 213;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 214;
address_inb = 215;
data_ina = 16'hfffe;
data_inb = 16'h1;
#10;
address_ina = 216;
address_inb = 217;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 218;
address_inb = 219;
data_ina = 16'hffff;
data_inb = 16'hfffe;
#10;
address_ina = 220;
address_inb = 221;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 222;
address_inb = 223;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 224;
address_inb = 225;
data_ina = 16'h0;
data_inb = 16'hfffd;
#10;
address_ina = 226;
address_inb = 227;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 228;
address_inb = 229;
data_ina = 16'h0;
data_inb = 16'hfffe;
#10;
address_ina = 230;
address_inb = 231;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 232;
address_inb = 233;
data_ina = 16'h2;
data_inb = 16'hffff;
#10;
address_ina = 234;
address_inb = 235;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 236;
address_inb = 237;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 238;
address_inb = 239;
data_ina = 16'h2;
data_inb = 16'h1;
#10;
address_ina = 240;
address_inb = 241;
data_ina = 16'hfffe;
data_inb = 16'hffff;
#10;
address_ina = 242;
address_inb = 243;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 244;
address_inb = 245;
data_ina = 16'h1;
data_inb = 16'hfffd;
#10;
address_ina = 246;
address_inb = 247;
data_ina = 16'h2;
data_inb = 16'h1;
#10;
address_ina = 248;
address_inb = 249;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 250;
address_inb = 251;
data_ina = 16'h1;
data_inb = 16'h3;
#10;
address_ina = 252;
address_inb = 253;
data_ina = 16'h0;
data_inb = 16'hfffd;
#10;
address_ina = 254;
address_inb = 255;
data_ina = 16'h1;
data_inb = 16'hfffe;
#10;
        wait(init_done);
        #30
        we = 0;
        // Start processing
         
		  #38000

        start = 0;



//        wait (wr_req);
//		  wait (!wr_req);
//		   rd_req = 1;
		  wait(done);
		  #20000
rd_req = 1;
        #70 
		  start = 1;
		 #80 
wait(rd_empty)
rd_req = 0;

$display("Finished the NTT test Number %d",test_num);
////Begin test number #55//////////////
rst = 1;

//#1000
start = 1;
mode = 0; //NTT 0 // INTT 1

// Reset for a few clock cycles

#1000

rst = 0;
test_num = test_num + 1;
#1000
we = 1;
address_ina = 0;
address_inb = 1;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 2;
address_inb = 3;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 4;
address_inb = 5;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 6;
address_inb = 7;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 8;
address_inb = 9;
data_ina = 16'h2;
data_inb = 16'h0;
#10;
address_ina = 10;
address_inb = 11;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 12;
address_inb = 13;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 14;
address_inb = 15;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 16;
address_inb = 17;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 18;
address_inb = 19;
data_ina = 16'hfffd;
data_inb = 16'h1;
#10;
address_ina = 20;
address_inb = 21;
data_ina = 16'h1;
data_inb = 16'h2;
#10;
address_ina = 22;
address_inb = 23;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 24;
address_inb = 25;
data_ina = 16'h1;
data_inb = 16'h2;
#10;
address_ina = 26;
address_inb = 27;
data_ina = 16'h2;
data_inb = 16'h1;
#10;
address_ina = 28;
address_inb = 29;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 30;
address_inb = 31;
data_ina = 16'h2;
data_inb = 16'h2;
#10;
address_ina = 32;
address_inb = 33;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 34;
address_inb = 35;
data_ina = 16'h0;
data_inb = 16'hfffe;
#10;
address_ina = 36;
address_inb = 37;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 38;
address_inb = 39;
data_ina = 16'hfffe;
data_inb = 16'hffff;
#10;
address_ina = 40;
address_inb = 41;
data_ina = 16'h0;
data_inb = 16'hfffd;
#10;
address_ina = 42;
address_inb = 43;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 44;
address_inb = 45;
data_ina = 16'hfffe;
data_inb = 16'hffff;
#10;
address_ina = 46;
address_inb = 47;
data_ina = 16'h3;
data_inb = 16'hfffd;
#10;
address_ina = 48;
address_inb = 49;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 50;
address_inb = 51;
data_ina = 16'h3;
data_inb = 16'h0;
#10;
address_ina = 52;
address_inb = 53;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 54;
address_inb = 55;
data_ina = 16'hfffd;
data_inb = 16'h1;
#10;
address_ina = 56;
address_inb = 57;
data_ina = 16'hffff;
data_inb = 16'hfffe;
#10;
address_ina = 58;
address_inb = 59;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 60;
address_inb = 61;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 62;
address_inb = 63;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 64;
address_inb = 65;
data_ina = 16'hfffe;
data_inb = 16'h1;
#10;
address_ina = 66;
address_inb = 67;
data_ina = 16'h2;
data_inb = 16'h2;
#10;
address_ina = 68;
address_inb = 69;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 70;
address_inb = 71;
data_ina = 16'hfffe;
data_inb = 16'hfffd;
#10;
address_ina = 72;
address_inb = 73;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 74;
address_inb = 75;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 76;
address_inb = 77;
data_ina = 16'hffff;
data_inb = 16'h2;
#10;
address_ina = 78;
address_inb = 79;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 80;
address_inb = 81;
data_ina = 16'h0;
data_inb = 16'hfffe;
#10;
address_ina = 82;
address_inb = 83;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 84;
address_inb = 85;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 86;
address_inb = 87;
data_ina = 16'h2;
data_inb = 16'h0;
#10;
address_ina = 88;
address_inb = 89;
data_ina = 16'h3;
data_inb = 16'hffff;
#10;
address_ina = 90;
address_inb = 91;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 92;
address_inb = 93;
data_ina = 16'hffff;
data_inb = 16'hfffd;
#10;
address_ina = 94;
address_inb = 95;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 96;
address_inb = 97;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 98;
address_inb = 99;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 100;
address_inb = 101;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 102;
address_inb = 103;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 104;
address_inb = 105;
data_ina = 16'h2;
data_inb = 16'h1;
#10;
address_ina = 106;
address_inb = 107;
data_ina = 16'hffff;
data_inb = 16'h2;
#10;
address_ina = 108;
address_inb = 109;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 110;
address_inb = 111;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 112;
address_inb = 113;
data_ina = 16'h0;
data_inb = 16'h3;
#10;
address_ina = 114;
address_inb = 115;
data_ina = 16'hfffe;
data_inb = 16'h1;
#10;
address_ina = 116;
address_inb = 117;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 118;
address_inb = 119;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 120;
address_inb = 121;
data_ina = 16'hfffe;
data_inb = 16'hfffe;
#10;
address_ina = 122;
address_inb = 123;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 124;
address_inb = 125;
data_ina = 16'h0;
data_inb = 16'hfffe;
#10;
address_ina = 126;
address_inb = 127;
data_ina = 16'h2;
data_inb = 16'hfffe;
#10;
address_ina = 128;
address_inb = 129;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 130;
address_inb = 131;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 132;
address_inb = 133;
data_ina = 16'hffff;
data_inb = 16'hfffe;
#10;
address_ina = 134;
address_inb = 135;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 136;
address_inb = 137;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 138;
address_inb = 139;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 140;
address_inb = 141;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 142;
address_inb = 143;
data_ina = 16'h2;
data_inb = 16'h1;
#10;
address_ina = 144;
address_inb = 145;
data_ina = 16'hffff;
data_inb = 16'hfffe;
#10;
address_ina = 146;
address_inb = 147;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 148;
address_inb = 149;
data_ina = 16'h0;
data_inb = 16'hfffe;
#10;
address_ina = 150;
address_inb = 151;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 152;
address_inb = 153;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 154;
address_inb = 155;
data_ina = 16'hfffd;
data_inb = 16'h1;
#10;
address_ina = 156;
address_inb = 157;
data_ina = 16'h2;
data_inb = 16'hffff;
#10;
address_ina = 158;
address_inb = 159;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 160;
address_inb = 161;
data_ina = 16'h3;
data_inb = 16'h0;
#10;
address_ina = 162;
address_inb = 163;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 164;
address_inb = 165;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 166;
address_inb = 167;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 168;
address_inb = 169;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 170;
address_inb = 171;
data_ina = 16'h1;
data_inb = 16'h3;
#10;
address_ina = 172;
address_inb = 173;
data_ina = 16'h0;
data_inb = 16'h2;
#10;
address_ina = 174;
address_inb = 175;
data_ina = 16'h1;
data_inb = 16'h3;
#10;
address_ina = 176;
address_inb = 177;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 178;
address_inb = 179;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 180;
address_inb = 181;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 182;
address_inb = 183;
data_ina = 16'hfffd;
data_inb = 16'h0;
#10;
address_ina = 184;
address_inb = 185;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 186;
address_inb = 187;
data_ina = 16'h3;
data_inb = 16'hffff;
#10;
address_ina = 188;
address_inb = 189;
data_ina = 16'hffff;
data_inb = 16'hfffe;
#10;
address_ina = 190;
address_inb = 191;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 192;
address_inb = 193;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 194;
address_inb = 195;
data_ina = 16'h2;
data_inb = 16'h0;
#10;
address_ina = 196;
address_inb = 197;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 198;
address_inb = 199;
data_ina = 16'h0;
data_inb = 16'h2;
#10;
address_ina = 200;
address_inb = 201;
data_ina = 16'hfffe;
data_inb = 16'h0;
#10;
address_ina = 202;
address_inb = 203;
data_ina = 16'h2;
data_inb = 16'h0;
#10;
address_ina = 204;
address_inb = 205;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 206;
address_inb = 207;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 208;
address_inb = 209;
data_ina = 16'h1;
data_inb = 16'h2;
#10;
address_ina = 210;
address_inb = 211;
data_ina = 16'hffff;
data_inb = 16'h2;
#10;
address_ina = 212;
address_inb = 213;
data_ina = 16'hfffe;
data_inb = 16'h1;
#10;
address_ina = 214;
address_inb = 215;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 216;
address_inb = 217;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 218;
address_inb = 219;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 220;
address_inb = 221;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 222;
address_inb = 223;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 224;
address_inb = 225;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 226;
address_inb = 227;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 228;
address_inb = 229;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 230;
address_inb = 231;
data_ina = 16'h1;
data_inb = 16'hfffd;
#10;
address_ina = 232;
address_inb = 233;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 234;
address_inb = 235;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 236;
address_inb = 237;
data_ina = 16'hfffe;
data_inb = 16'h1;
#10;
address_ina = 238;
address_inb = 239;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 240;
address_inb = 241;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 242;
address_inb = 243;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 244;
address_inb = 245;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 246;
address_inb = 247;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 248;
address_inb = 249;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 250;
address_inb = 251;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 252;
address_inb = 253;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 254;
address_inb = 255;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
        wait(init_done);
        #30
        we = 0;
        // Start processing
         
		  #38000

        start = 0;



//        wait (wr_req);
//		  wait (!wr_req);
//		   rd_req = 1;
		  wait(done);
		  #20000
rd_req = 1;
        #70 
		  start = 1;
		 #80 
wait(rd_empty)
rd_req = 0;

$display("Finished the NTT test Number %d",test_num);
////Begin test number #56//////////////
rst = 1;

//#1000
start = 1;
mode = 0; //NTT 0 // INTT 1

// Reset for a few clock cycles

#1000

rst = 0;
test_num = test_num + 1;
#1000
we = 1;
address_ina = 0;
address_inb = 1;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 2;
address_inb = 3;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 4;
address_inb = 5;
data_ina = 16'hfffe;
data_inb = 16'h1;
#10;
address_ina = 6;
address_inb = 7;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 8;
address_inb = 9;
data_ina = 16'h3;
data_inb = 16'h0;
#10;
address_ina = 10;
address_inb = 11;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 12;
address_inb = 13;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 14;
address_inb = 15;
data_ina = 16'hffff;
data_inb = 16'hfffe;
#10;
address_ina = 16;
address_inb = 17;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 18;
address_inb = 19;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 20;
address_inb = 21;
data_ina = 16'hfffe;
data_inb = 16'h0;
#10;
address_ina = 22;
address_inb = 23;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 24;
address_inb = 25;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 26;
address_inb = 27;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 28;
address_inb = 29;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 30;
address_inb = 31;
data_ina = 16'h1;
data_inb = 16'h3;
#10;
address_ina = 32;
address_inb = 33;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 34;
address_inb = 35;
data_ina = 16'hfffe;
data_inb = 16'h1;
#10;
address_ina = 36;
address_inb = 37;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 38;
address_inb = 39;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 40;
address_inb = 41;
data_ina = 16'h0;
data_inb = 16'hfffe;
#10;
address_ina = 42;
address_inb = 43;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 44;
address_inb = 45;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 46;
address_inb = 47;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 48;
address_inb = 49;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 50;
address_inb = 51;
data_ina = 16'hfffe;
data_inb = 16'hffff;
#10;
address_ina = 52;
address_inb = 53;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 54;
address_inb = 55;
data_ina = 16'h1;
data_inb = 16'hfffd;
#10;
address_ina = 56;
address_inb = 57;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 58;
address_inb = 59;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 60;
address_inb = 61;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 62;
address_inb = 63;
data_ina = 16'hfffe;
data_inb = 16'h0;
#10;
address_ina = 64;
address_inb = 65;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 66;
address_inb = 67;
data_ina = 16'hffff;
data_inb = 16'hfffe;
#10;
address_ina = 68;
address_inb = 69;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 70;
address_inb = 71;
data_ina = 16'h0;
data_inb = 16'h2;
#10;
address_ina = 72;
address_inb = 73;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 74;
address_inb = 75;
data_ina = 16'h1;
data_inb = 16'hfffe;
#10;
address_ina = 76;
address_inb = 77;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 78;
address_inb = 79;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 80;
address_inb = 81;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 82;
address_inb = 83;
data_ina = 16'hffff;
data_inb = 16'h2;
#10;
address_ina = 84;
address_inb = 85;
data_ina = 16'h2;
data_inb = 16'hfffd;
#10;
address_ina = 86;
address_inb = 87;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 88;
address_inb = 89;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 90;
address_inb = 91;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 92;
address_inb = 93;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 94;
address_inb = 95;
data_ina = 16'h1;
data_inb = 16'hfffe;
#10;
address_ina = 96;
address_inb = 97;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 98;
address_inb = 99;
data_ina = 16'h0;
data_inb = 16'h2;
#10;
address_ina = 100;
address_inb = 101;
data_ina = 16'hfffe;
data_inb = 16'hffff;
#10;
address_ina = 102;
address_inb = 103;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 104;
address_inb = 105;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 106;
address_inb = 107;
data_ina = 16'h2;
data_inb = 16'hffff;
#10;
address_ina = 108;
address_inb = 109;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 110;
address_inb = 111;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 112;
address_inb = 113;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 114;
address_inb = 115;
data_ina = 16'h2;
data_inb = 16'h1;
#10;
address_ina = 116;
address_inb = 117;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 118;
address_inb = 119;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 120;
address_inb = 121;
data_ina = 16'hfffe;
data_inb = 16'h1;
#10;
address_ina = 122;
address_inb = 123;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 124;
address_inb = 125;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 126;
address_inb = 127;
data_ina = 16'h2;
data_inb = 16'h0;
#10;
address_ina = 128;
address_inb = 129;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 130;
address_inb = 131;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 132;
address_inb = 133;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 134;
address_inb = 135;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 136;
address_inb = 137;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 138;
address_inb = 139;
data_ina = 16'hffff;
data_inb = 16'h2;
#10;
address_ina = 140;
address_inb = 141;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 142;
address_inb = 143;
data_ina = 16'h1;
data_inb = 16'hfffe;
#10;
address_ina = 144;
address_inb = 145;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 146;
address_inb = 147;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 148;
address_inb = 149;
data_ina = 16'h2;
data_inb = 16'h2;
#10;
address_ina = 150;
address_inb = 151;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 152;
address_inb = 153;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 154;
address_inb = 155;
data_ina = 16'hffff;
data_inb = 16'h2;
#10;
address_ina = 156;
address_inb = 157;
data_ina = 16'hfffe;
data_inb = 16'hffff;
#10;
address_ina = 158;
address_inb = 159;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 160;
address_inb = 161;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 162;
address_inb = 163;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 164;
address_inb = 165;
data_ina = 16'hfffd;
data_inb = 16'hffff;
#10;
address_ina = 166;
address_inb = 167;
data_ina = 16'hfffe;
data_inb = 16'h0;
#10;
address_ina = 168;
address_inb = 169;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 170;
address_inb = 171;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 172;
address_inb = 173;
data_ina = 16'h1;
data_inb = 16'hfffe;
#10;
address_ina = 174;
address_inb = 175;
data_ina = 16'hfffe;
data_inb = 16'h1;
#10;
address_ina = 176;
address_inb = 177;
data_ina = 16'hffff;
data_inb = 16'h2;
#10;
address_ina = 178;
address_inb = 179;
data_ina = 16'hfffe;
data_inb = 16'h0;
#10;
address_ina = 180;
address_inb = 181;
data_ina = 16'h1;
data_inb = 16'h2;
#10;
address_ina = 182;
address_inb = 183;
data_ina = 16'hffff;
data_inb = 16'h3;
#10;
address_ina = 184;
address_inb = 185;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 186;
address_inb = 187;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 188;
address_inb = 189;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 190;
address_inb = 191;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 192;
address_inb = 193;
data_ina = 16'hffff;
data_inb = 16'hfffe;
#10;
address_ina = 194;
address_inb = 195;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 196;
address_inb = 197;
data_ina = 16'h0;
data_inb = 16'hfffe;
#10;
address_ina = 198;
address_inb = 199;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 200;
address_inb = 201;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 202;
address_inb = 203;
data_ina = 16'h2;
data_inb = 16'h0;
#10;
address_ina = 204;
address_inb = 205;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 206;
address_inb = 207;
data_ina = 16'hfffd;
data_inb = 16'hfffe;
#10;
address_ina = 208;
address_inb = 209;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 210;
address_inb = 211;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 212;
address_inb = 213;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 214;
address_inb = 215;
data_ina = 16'h0;
data_inb = 16'h2;
#10;
address_ina = 216;
address_inb = 217;
data_ina = 16'h2;
data_inb = 16'h1;
#10;
address_ina = 218;
address_inb = 219;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 220;
address_inb = 221;
data_ina = 16'h3;
data_inb = 16'h1;
#10;
address_ina = 222;
address_inb = 223;
data_ina = 16'h2;
data_inb = 16'hffff;
#10;
address_ina = 224;
address_inb = 225;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 226;
address_inb = 227;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 228;
address_inb = 229;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 230;
address_inb = 231;
data_ina = 16'h2;
data_inb = 16'h1;
#10;
address_ina = 232;
address_inb = 233;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 234;
address_inb = 235;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 236;
address_inb = 237;
data_ina = 16'h0;
data_inb = 16'hfffe;
#10;
address_ina = 238;
address_inb = 239;
data_ina = 16'h0;
data_inb = 16'hfffe;
#10;
address_ina = 240;
address_inb = 241;
data_ina = 16'hfffe;
data_inb = 16'hfffe;
#10;
address_ina = 242;
address_inb = 243;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 244;
address_inb = 245;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 246;
address_inb = 247;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 248;
address_inb = 249;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 250;
address_inb = 251;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 252;
address_inb = 253;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 254;
address_inb = 255;
data_ina = 16'h1;
data_inb = 16'h2;
#10;
        wait(init_done);
        #30
        we = 0;
        // Start processing
         
		  #38000

        start = 0;



//        wait (wr_req);
//		  wait (!wr_req);
//		   rd_req = 1;
		  wait(done);
		  #20000
rd_req = 1;
        #70 
		  start = 1;
		 #80 
wait(rd_empty)
rd_req = 0;

$display("Finished the NTT test Number %d",test_num);
////Begin test number #57//////////////
rst = 1;

//#1000
start = 1;
mode = 1; //NTT 0 // INTT 1

// Reset for a few clock cycles

#1000

rst = 0;
test_num = test_num + 1;
#1000
we = 1;
address_ina = 0;
address_inb = 1;
data_ina = 16'hfc36;
data_inb = 16'ha5;
#10;
address_ina = 2;
address_inb = 3;
data_ina = 16'h4b3;
data_inb = 16'h22b;
#10;
address_ina = 4;
address_inb = 5;
data_ina = 16'hfb68;
data_inb = 16'hc4;
#10;
address_ina = 6;
address_inb = 7;
data_ina = 16'hfb62;
data_inb = 16'hfb88;
#10;
address_ina = 8;
address_inb = 9;
data_ina = 16'hf0;
data_inb = 16'hfa50;
#10;
address_ina = 10;
address_inb = 11;
data_ina = 16'hfb45;
data_inb = 16'h17;
#10;
address_ina = 12;
address_inb = 13;
data_ina = 16'h11c;
data_inb = 16'hc0;
#10;
address_ina = 14;
address_inb = 15;
data_ina = 16'hfa7e;
data_inb = 16'hfdd0;
#10;
address_ina = 16;
address_inb = 17;
data_ina = 16'hff51;
data_inb = 16'h468;
#10;
address_ina = 18;
address_inb = 19;
data_ina = 16'hfd2a;
data_inb = 16'h30b;
#10;
address_ina = 20;
address_inb = 21;
data_ina = 16'h412;
data_inb = 16'hfeb3;
#10;
address_ina = 22;
address_inb = 23;
data_ina = 16'h50b;
data_inb = 16'hfbe6;
#10;
address_ina = 24;
address_inb = 25;
data_ina = 16'hfb43;
data_inb = 16'h3ee;
#10;
address_ina = 26;
address_inb = 27;
data_ina = 16'h196;
data_inb = 16'hff28;
#10;
address_ina = 28;
address_inb = 29;
data_ina = 16'hfe59;
data_inb = 16'hfa6d;
#10;
address_ina = 30;
address_inb = 31;
data_ina = 16'h3b5;
data_inb = 16'h593;
#10;
address_ina = 32;
address_inb = 33;
data_ina = 16'hfb2e;
data_inb = 16'hfeb4;
#10;
address_ina = 34;
address_inb = 35;
data_ina = 16'h475;
data_inb = 16'h386;
#10;
address_ina = 36;
address_inb = 37;
data_ina = 16'hfab1;
data_inb = 16'h3f4;
#10;
address_ina = 38;
address_inb = 39;
data_ina = 16'hfe17;
data_inb = 16'hfc5e;
#10;
address_ina = 40;
address_inb = 41;
data_ina = 16'hfe8c;
data_inb = 16'hfcd6;
#10;
address_ina = 42;
address_inb = 43;
data_ina = 16'hfa34;
data_inb = 16'hfbc8;
#10;
address_ina = 44;
address_inb = 45;
data_ina = 16'h3d9;
data_inb = 16'h40b;
#10;
address_ina = 46;
address_inb = 47;
data_ina = 16'hf9ed;
data_inb = 16'h32;
#10;
address_ina = 48;
address_inb = 49;
data_ina = 16'h282;
data_inb = 16'h52;
#10;
address_ina = 50;
address_inb = 51;
data_ina = 16'hf9c5;
data_inb = 16'h4bb;
#10;
address_ina = 52;
address_inb = 53;
data_ina = 16'hfd1d;
data_inb = 16'h7a;
#10;
address_ina = 54;
address_inb = 55;
data_ina = 16'hfa8e;
data_inb = 16'hff38;
#10;
address_ina = 56;
address_inb = 57;
data_ina = 16'h22;
data_inb = 16'hfc59;
#10;
address_ina = 58;
address_inb = 59;
data_ina = 16'h51c;
data_inb = 16'h581;
#10;
address_ina = 60;
address_inb = 61;
data_ina = 16'hfb57;
data_inb = 16'h542;
#10;
address_ina = 62;
address_inb = 63;
data_ina = 16'h608;
data_inb = 16'h573;
#10;
address_ina = 64;
address_inb = 65;
data_ina = 16'h535;
data_inb = 16'hff9e;
#10;
address_ina = 66;
address_inb = 67;
data_ina = 16'hfe9a;
data_inb = 16'hfa3d;
#10;
address_ina = 68;
address_inb = 69;
data_ina = 16'h2a;
data_inb = 16'h671;
#10;
address_ina = 70;
address_inb = 71;
data_ina = 16'hffc4;
data_inb = 16'h59a;
#10;
address_ina = 72;
address_inb = 73;
data_ina = 16'hfb05;
data_inb = 16'hf995;
#10;
address_ina = 74;
address_inb = 75;
data_ina = 16'h352;
data_inb = 16'hfc88;
#10;
address_ina = 76;
address_inb = 77;
data_ina = 16'h642;
data_inb = 16'hfd4c;
#10;
address_ina = 78;
address_inb = 79;
data_ina = 16'hfdea;
data_inb = 16'hffb2;
#10;
address_ina = 80;
address_inb = 81;
data_ina = 16'hfb18;
data_inb = 16'hfd53;
#10;
address_ina = 82;
address_inb = 83;
data_ina = 16'hfaf7;
data_inb = 16'h5f6;
#10;
address_ina = 84;
address_inb = 85;
data_ina = 16'h67a;
data_inb = 16'hff9c;
#10;
address_ina = 86;
address_inb = 87;
data_ina = 16'h566;
data_inb = 16'h302;
#10;
address_ina = 88;
address_inb = 89;
data_ina = 16'h2fa;
data_inb = 16'h4e2;
#10;
address_ina = 90;
address_inb = 91;
data_ina = 16'h411;
data_inb = 16'hfbe2;
#10;
address_ina = 92;
address_inb = 93;
data_ina = 16'hfe68;
data_inb = 16'hf9a7;
#10;
address_ina = 94;
address_inb = 95;
data_ina = 16'hfd7b;
data_inb = 16'h32b;
#10;
address_ina = 96;
address_inb = 97;
data_ina = 16'h7f;
data_inb = 16'hfdbc;
#10;
address_ina = 98;
address_inb = 99;
data_ina = 16'hfc59;
data_inb = 16'hfb21;
#10;
address_ina = 100;
address_inb = 101;
data_ina = 16'hff3c;
data_inb = 16'h2a7;
#10;
address_ina = 102;
address_inb = 103;
data_ina = 16'h3f2;
data_inb = 16'h623;
#10;
address_ina = 104;
address_inb = 105;
data_ina = 16'h56e;
data_inb = 16'hfe29;
#10;
address_ina = 106;
address_inb = 107;
data_ina = 16'h57;
data_inb = 16'hfd15;
#10;
address_ina = 108;
address_inb = 109;
data_ina = 16'hfee6;
data_inb = 16'hff88;
#10;
address_ina = 110;
address_inb = 111;
data_ina = 16'h518;
data_inb = 16'h627;
#10;
address_ina = 112;
address_inb = 113;
data_ina = 16'h435;
data_inb = 16'h302;
#10;
address_ina = 114;
address_inb = 115;
data_ina = 16'hfb00;
data_inb = 16'h298;
#10;
address_ina = 116;
address_inb = 117;
data_ina = 16'hfb3f;
data_inb = 16'hf9eb;
#10;
address_ina = 118;
address_inb = 119;
data_ina = 16'h623;
data_inb = 16'hfb86;
#10;
address_ina = 120;
address_inb = 121;
data_ina = 16'hf9dc;
data_inb = 16'hf997;
#10;
address_ina = 122;
address_inb = 123;
data_ina = 16'hfacf;
data_inb = 16'hffef;
#10;
address_ina = 124;
address_inb = 125;
data_ina = 16'hfe6f;
data_inb = 16'h1e5;
#10;
address_ina = 126;
address_inb = 127;
data_ina = 16'h52a;
data_inb = 16'hfbc0;
#10;
address_ina = 128;
address_inb = 129;
data_ina = 16'h89;
data_inb = 16'h455;
#10;
address_ina = 130;
address_inb = 131;
data_ina = 16'hfa22;
data_inb = 16'hff5b;
#10;
address_ina = 132;
address_inb = 133;
data_ina = 16'h269;
data_inb = 16'hfce6;
#10;
address_ina = 134;
address_inb = 135;
data_ina = 16'hff5e;
data_inb = 16'hfd1c;
#10;
address_ina = 136;
address_inb = 137;
data_ina = 16'hfedd;
data_inb = 16'hffae;
#10;
address_ina = 138;
address_inb = 139;
data_ina = 16'h667;
data_inb = 16'h3a3;
#10;
address_ina = 140;
address_inb = 141;
data_ina = 16'h4dd;
data_inb = 16'h16f;
#10;
address_ina = 142;
address_inb = 143;
data_ina = 16'h535;
data_inb = 16'h344;
#10;
address_ina = 144;
address_inb = 145;
data_ina = 16'hff25;
data_inb = 16'h159;
#10;
address_ina = 146;
address_inb = 147;
data_ina = 16'hf9b7;
data_inb = 16'hfe91;
#10;
address_ina = 148;
address_inb = 149;
data_ina = 16'h4aa;
data_inb = 16'hfa15;
#10;
address_ina = 150;
address_inb = 151;
data_ina = 16'hfa82;
data_inb = 16'h536;
#10;
address_ina = 152;
address_inb = 153;
data_ina = 16'hffe7;
data_inb = 16'h3b2;
#10;
address_ina = 154;
address_inb = 155;
data_ina = 16'h85;
data_inb = 16'h183;
#10;
address_ina = 156;
address_inb = 157;
data_ina = 16'hfa43;
data_inb = 16'h242;
#10;
address_ina = 158;
address_inb = 159;
data_ina = 16'hfc4a;
data_inb = 16'hfb26;
#10;
address_ina = 160;
address_inb = 161;
data_ina = 16'hfec8;
data_inb = 16'hfc3b;
#10;
address_ina = 162;
address_inb = 163;
data_ina = 16'h303;
data_inb = 16'hff37;
#10;
address_ina = 164;
address_inb = 165;
data_ina = 16'h50;
data_inb = 16'hf9b8;
#10;
address_ina = 166;
address_inb = 167;
data_ina = 16'h633;
data_inb = 16'hfe11;
#10;
address_ina = 168;
address_inb = 169;
data_ina = 16'hff1e;
data_inb = 16'hfc48;
#10;
address_ina = 170;
address_inb = 171;
data_ina = 16'hfa1c;
data_inb = 16'hf9c6;
#10;
address_ina = 172;
address_inb = 173;
data_ina = 16'h5f3;
data_inb = 16'h666;
#10;
address_ina = 174;
address_inb = 175;
data_ina = 16'h15e;
data_inb = 16'h1a5;
#10;
address_ina = 176;
address_inb = 177;
data_ina = 16'hfed5;
data_inb = 16'hfbfd;
#10;
address_ina = 178;
address_inb = 179;
data_ina = 16'h5fd;
data_inb = 16'h507;
#10;
address_ina = 180;
address_inb = 181;
data_ina = 16'hfa83;
data_inb = 16'hff18;
#10;
address_ina = 182;
address_inb = 183;
data_ina = 16'h9;
data_inb = 16'hfcba;
#10;
address_ina = 184;
address_inb = 185;
data_ina = 16'h290;
data_inb = 16'hfce8;
#10;
address_ina = 186;
address_inb = 187;
data_ina = 16'hfb2f;
data_inb = 16'hfdac;
#10;
address_ina = 188;
address_inb = 189;
data_ina = 16'hfd68;
data_inb = 16'hfea9;
#10;
address_ina = 190;
address_inb = 191;
data_ina = 16'h3c7;
data_inb = 16'h45a;
#10;
address_ina = 192;
address_inb = 193;
data_ina = 16'hfc4d;
data_inb = 16'hfa8a;
#10;
address_ina = 194;
address_inb = 195;
data_ina = 16'h2ad;
data_inb = 16'hfcfe;
#10;
address_ina = 196;
address_inb = 197;
data_ina = 16'h33f;
data_inb = 16'hfb04;
#10;
address_ina = 198;
address_inb = 199;
data_ina = 16'hfeaf;
data_inb = 16'hfa3d;
#10;
address_ina = 200;
address_inb = 201;
data_ina = 16'h601;
data_inb = 16'h3cb;
#10;
address_ina = 202;
address_inb = 203;
data_ina = 16'h40c;
data_inb = 16'h67;
#10;
address_ina = 204;
address_inb = 205;
data_ina = 16'hfbf0;
data_inb = 16'hb7;
#10;
address_ina = 206;
address_inb = 207;
data_ina = 16'hff8b;
data_inb = 16'hfc6b;
#10;
address_ina = 208;
address_inb = 209;
data_ina = 16'h396;
data_inb = 16'h363;
#10;
address_ina = 210;
address_inb = 211;
data_ina = 16'hfc53;
data_inb = 16'hff01;
#10;
address_ina = 212;
address_inb = 213;
data_ina = 16'hfee7;
data_inb = 16'h190;
#10;
address_ina = 214;
address_inb = 215;
data_ina = 16'h492;
data_inb = 16'h8b;
#10;
address_ina = 216;
address_inb = 217;
data_ina = 16'hff9b;
data_inb = 16'hfdfd;
#10;
address_ina = 218;
address_inb = 219;
data_ina = 16'he7;
data_inb = 16'h675;
#10;
address_ina = 220;
address_inb = 221;
data_ina = 16'h24a;
data_inb = 16'h26a;
#10;
address_ina = 222;
address_inb = 223;
data_ina = 16'h4fd;
data_inb = 16'h284;
#10;
address_ina = 224;
address_inb = 225;
data_ina = 16'hfab6;
data_inb = 16'hfc5f;
#10;
address_ina = 226;
address_inb = 227;
data_ina = 16'hfc6b;
data_inb = 16'h4fe;
#10;
address_ina = 228;
address_inb = 229;
data_ina = 16'h295;
data_inb = 16'hfe96;
#10;
address_ina = 230;
address_inb = 231;
data_ina = 16'hfb96;
data_inb = 16'hfeac;
#10;
address_ina = 232;
address_inb = 233;
data_ina = 16'hf4;
data_inb = 16'h9d;
#10;
address_ina = 234;
address_inb = 235;
data_ina = 16'hfb27;
data_inb = 16'hfd89;
#10;
address_ina = 236;
address_inb = 237;
data_ina = 16'h1b3;
data_inb = 16'hd9;
#10;
address_ina = 238;
address_inb = 239;
data_ina = 16'h171;
data_inb = 16'hfb45;
#10;
address_ina = 240;
address_inb = 241;
data_ina = 16'hfffb;
data_inb = 16'hf985;
#10;
address_ina = 242;
address_inb = 243;
data_ina = 16'h400;
data_inb = 16'hfc81;
#10;
address_ina = 244;
address_inb = 245;
data_ina = 16'hfd6f;
data_inb = 16'h39a;
#10;
address_ina = 246;
address_inb = 247;
data_ina = 16'h4dd;
data_inb = 16'hfb0b;
#10;
address_ina = 248;
address_inb = 249;
data_ina = 16'hfaad;
data_inb = 16'hf9ab;
#10;
address_ina = 250;
address_inb = 251;
data_ina = 16'h599;
data_inb = 16'h44f;
#10;
address_ina = 252;
address_inb = 253;
data_ina = 16'h4dc;
data_inb = 16'hfc75;
#10;
address_ina = 254;
address_inb = 255;
data_ina = 16'h59c;
data_inb = 16'h1ec;
#10;
        wait(init_done);
        #30
        we = 0;
        // Start processing
         
		  #38000

        start = 0;



//        wait (wr_req);
//		  wait (!wr_req);
//		   rd_req = 1;
		  wait(done);
		  #20000
rd_req = 1;
        #70 
		  start = 1;
		 #80 
wait(rd_empty)
rd_req = 0;

$display("Finished the NTT test Number %d",test_num);
////Begin test number #58//////////////
rst = 1;

//#1000
start = 1;
mode = 1; //NTT 0 // INTT 1

// Reset for a few clock cycles

#1000

rst = 0;
test_num = test_num + 1;
#1000
we = 1;
address_ina = 0;
address_inb = 1;
data_ina = 16'hfd7b;
data_inb = 16'hfd91;
#10;
address_ina = 2;
address_inb = 3;
data_ina = 16'h5da;
data_inb = 16'h24c;
#10;
address_ina = 4;
address_inb = 5;
data_ina = 16'h59b;
data_inb = 16'h64a;
#10;
address_ina = 6;
address_inb = 7;
data_ina = 16'h594;
data_inb = 16'hfad7;
#10;
address_ina = 8;
address_inb = 9;
data_ina = 16'hf993;
data_inb = 16'h2b2;
#10;
address_ina = 10;
address_inb = 11;
data_ina = 16'ha;
data_inb = 16'hffcc;
#10;
address_ina = 12;
address_inb = 13;
data_ina = 16'hfeb7;
data_inb = 16'hf9d8;
#10;
address_ina = 14;
address_inb = 15;
data_ina = 16'h3ae;
data_inb = 16'hfd50;
#10;
address_ina = 16;
address_inb = 17;
data_ina = 16'h550;
data_inb = 16'hf9a2;
#10;
address_ina = 18;
address_inb = 19;
data_ina = 16'hfceb;
data_inb = 16'h567;
#10;
address_ina = 20;
address_inb = 21;
data_ina = 16'h121;
data_inb = 16'h182;
#10;
address_ina = 22;
address_inb = 23;
data_ina = 16'h65f;
data_inb = 16'h4bf;
#10;
address_ina = 24;
address_inb = 25;
data_ina = 16'h135;
data_inb = 16'hde;
#10;
address_ina = 26;
address_inb = 27;
data_ina = 16'hfd7b;
data_inb = 16'h272;
#10;
address_ina = 28;
address_inb = 29;
data_ina = 16'h4ae;
data_inb = 16'h2ff;
#10;
address_ina = 30;
address_inb = 31;
data_ina = 16'hfa78;
data_inb = 16'h329;
#10;
address_ina = 32;
address_inb = 33;
data_ina = 16'hfc08;
data_inb = 16'h2ad;
#10;
address_ina = 34;
address_inb = 35;
data_ina = 16'hfa77;
data_inb = 16'hffbb;
#10;
address_ina = 36;
address_inb = 37;
data_ina = 16'hfe09;
data_inb = 16'hfb4d;
#10;
address_ina = 38;
address_inb = 39;
data_ina = 16'h502;
data_inb = 16'h1d6;
#10;
address_ina = 40;
address_inb = 41;
data_ina = 16'hfe48;
data_inb = 16'hffbd;
#10;
address_ina = 42;
address_inb = 43;
data_ina = 16'hfae6;
data_inb = 16'hfbbc;
#10;
address_ina = 44;
address_inb = 45;
data_ina = 16'h2ac;
data_inb = 16'h48c;
#10;
address_ina = 46;
address_inb = 47;
data_ina = 16'h3f6;
data_inb = 16'hfb3d;
#10;
address_ina = 48;
address_inb = 49;
data_ina = 16'hfbb3;
data_inb = 16'hfd24;
#10;
address_ina = 50;
address_inb = 51;
data_ina = 16'hfd44;
data_inb = 16'h318;
#10;
address_ina = 52;
address_inb = 53;
data_ina = 16'h44;
data_inb = 16'h660;
#10;
address_ina = 54;
address_inb = 55;
data_ina = 16'hfe6e;
data_inb = 16'hfe97;
#10;
address_ina = 56;
address_inb = 57;
data_ina = 16'hfe99;
data_inb = 16'h37c;
#10;
address_ina = 58;
address_inb = 59;
data_ina = 16'hfca0;
data_inb = 16'h593;
#10;
address_ina = 60;
address_inb = 61;
data_ina = 16'h283;
data_inb = 16'h1a5;
#10;
address_ina = 62;
address_inb = 63;
data_ina = 16'h80;
data_inb = 16'hfce0;
#10;
address_ina = 64;
address_inb = 65;
data_ina = 16'hf99e;
data_inb = 16'h53b;
#10;
address_ina = 66;
address_inb = 67;
data_ina = 16'h62d;
data_inb = 16'hff6f;
#10;
address_ina = 68;
address_inb = 69;
data_ina = 16'h408;
data_inb = 16'hff96;
#10;
address_ina = 70;
address_inb = 71;
data_ina = 16'h13f;
data_inb = 16'hfa23;
#10;
address_ina = 72;
address_inb = 73;
data_ina = 16'h1d6;
data_inb = 16'h53e;
#10;
address_ina = 74;
address_inb = 75;
data_ina = 16'hfd73;
data_inb = 16'hf989;
#10;
address_ina = 76;
address_inb = 77;
data_ina = 16'hfc97;
data_inb = 16'h241;
#10;
address_ina = 78;
address_inb = 79;
data_ina = 16'h375;
data_inb = 16'hff3e;
#10;
address_ina = 80;
address_inb = 81;
data_ina = 16'h574;
data_inb = 16'hfbd5;
#10;
address_ina = 82;
address_inb = 83;
data_ina = 16'h184;
data_inb = 16'h58f;
#10;
address_ina = 84;
address_inb = 85;
data_ina = 16'he7;
data_inb = 16'hfae1;
#10;
address_ina = 86;
address_inb = 87;
data_ina = 16'h137;
data_inb = 16'h1ad;
#10;
address_ina = 88;
address_inb = 89;
data_ina = 16'hfa13;
data_inb = 16'h15;
#10;
address_ina = 90;
address_inb = 91;
data_ina = 16'h48;
data_inb = 16'hfde1;
#10;
address_ina = 92;
address_inb = 93;
data_ina = 16'h203;
data_inb = 16'h3c7;
#10;
address_ina = 94;
address_inb = 95;
data_ina = 16'h433;
data_inb = 16'hfdff;
#10;
address_ina = 96;
address_inb = 97;
data_ina = 16'h545;
data_inb = 16'hfc5b;
#10;
address_ina = 98;
address_inb = 99;
data_ina = 16'hff9c;
data_inb = 16'h146;
#10;
address_ina = 100;
address_inb = 101;
data_ina = 16'h3a5;
data_inb = 16'hfdea;
#10;
address_ina = 102;
address_inb = 103;
data_ina = 16'h254;
data_inb = 16'h2a6;
#10;
address_ina = 104;
address_inb = 105;
data_ina = 16'hfba4;
data_inb = 16'h40;
#10;
address_ina = 106;
address_inb = 107;
data_ina = 16'h12;
data_inb = 16'h3a9;
#10;
address_ina = 108;
address_inb = 109;
data_ina = 16'h5fd;
data_inb = 16'h2e;
#10;
address_ina = 110;
address_inb = 111;
data_ina = 16'hfd58;
data_inb = 16'hffa6;
#10;
address_ina = 112;
address_inb = 113;
data_ina = 16'h424;
data_inb = 16'hfc4c;
#10;
address_ina = 114;
address_inb = 115;
data_ina = 16'h305;
data_inb = 16'h2bb;
#10;
address_ina = 116;
address_inb = 117;
data_ina = 16'h30a;
data_inb = 16'hfc37;
#10;
address_ina = 118;
address_inb = 119;
data_ina = 16'h13e;
data_inb = 16'h13;
#10;
address_ina = 120;
address_inb = 121;
data_ina = 16'h5e;
data_inb = 16'hfcc5;
#10;
address_ina = 122;
address_inb = 123;
data_ina = 16'h1c2;
data_inb = 16'hfd53;
#10;
address_ina = 124;
address_inb = 125;
data_ina = 16'hfb7e;
data_inb = 16'hfc93;
#10;
address_ina = 126;
address_inb = 127;
data_ina = 16'h5dc;
data_inb = 16'hfe89;
#10;
address_ina = 128;
address_inb = 129;
data_ina = 16'h2a1;
data_inb = 16'h153;
#10;
address_ina = 130;
address_inb = 131;
data_ina = 16'hfb2e;
data_inb = 16'hfb06;
#10;
address_ina = 132;
address_inb = 133;
data_ina = 16'hfe4e;
data_inb = 16'h252;
#10;
address_ina = 134;
address_inb = 135;
data_ina = 16'h55f;
data_inb = 16'h5ae;
#10;
address_ina = 136;
address_inb = 137;
data_ina = 16'h258;
data_inb = 16'hff8b;
#10;
address_ina = 138;
address_inb = 139;
data_ina = 16'h152;
data_inb = 16'hfe9d;
#10;
address_ina = 140;
address_inb = 141;
data_ina = 16'hfab3;
data_inb = 16'hfdb7;
#10;
address_ina = 142;
address_inb = 143;
data_ina = 16'h3b;
data_inb = 16'hfb3f;
#10;
address_ina = 144;
address_inb = 145;
data_ina = 16'h27b;
data_inb = 16'h432;
#10;
address_ina = 146;
address_inb = 147;
data_ina = 16'hfd47;
data_inb = 16'hfb61;
#10;
address_ina = 148;
address_inb = 149;
data_ina = 16'hfc9d;
data_inb = 16'h12a;
#10;
address_ina = 150;
address_inb = 151;
data_ina = 16'h5ec;
data_inb = 16'h313;
#10;
address_ina = 152;
address_inb = 153;
data_ina = 16'h639;
data_inb = 16'hfc0d;
#10;
address_ina = 154;
address_inb = 155;
data_ina = 16'hfcf5;
data_inb = 16'hfa88;
#10;
address_ina = 156;
address_inb = 157;
data_ina = 16'h340;
data_inb = 16'hfa63;
#10;
address_ina = 158;
address_inb = 159;
data_ina = 16'h596;
data_inb = 16'h5d9;
#10;
address_ina = 160;
address_inb = 161;
data_ina = 16'hfaa0;
data_inb = 16'hfb32;
#10;
address_ina = 162;
address_inb = 163;
data_ina = 16'h2ef;
data_inb = 16'hfece;
#10;
address_ina = 164;
address_inb = 165;
data_ina = 16'h23b;
data_inb = 16'h35a;
#10;
address_ina = 166;
address_inb = 167;
data_ina = 16'hfbfa;
data_inb = 16'h84;
#10;
address_ina = 168;
address_inb = 169;
data_ina = 16'h224;
data_inb = 16'h4bc;
#10;
address_ina = 170;
address_inb = 171;
data_ina = 16'h3a3;
data_inb = 16'hfe72;
#10;
address_ina = 172;
address_inb = 173;
data_ina = 16'hf9c5;
data_inb = 16'h50b;
#10;
address_ina = 174;
address_inb = 175;
data_ina = 16'h2cf;
data_inb = 16'hfaed;
#10;
address_ina = 176;
address_inb = 177;
data_ina = 16'h3e0;
data_inb = 16'h3a0;
#10;
address_ina = 178;
address_inb = 179;
data_ina = 16'h3cc;
data_inb = 16'hff3b;
#10;
address_ina = 180;
address_inb = 181;
data_ina = 16'h42c;
data_inb = 16'hfc14;
#10;
address_ina = 182;
address_inb = 183;
data_ina = 16'h5c1;
data_inb = 16'h524;
#10;
address_ina = 184;
address_inb = 185;
data_ina = 16'h36d;
data_inb = 16'h422;
#10;
address_ina = 186;
address_inb = 187;
data_ina = 16'h21a;
data_inb = 16'hfef0;
#10;
address_ina = 188;
address_inb = 189;
data_ina = 16'hfad8;
data_inb = 16'h219;
#10;
address_ina = 190;
address_inb = 191;
data_ina = 16'hfcb0;
data_inb = 16'h82;
#10;
address_ina = 192;
address_inb = 193;
data_ina = 16'hfd8e;
data_inb = 16'h2fd;
#10;
address_ina = 194;
address_inb = 195;
data_ina = 16'h104;
data_inb = 16'h120;
#10;
address_ina = 196;
address_inb = 197;
data_ina = 16'hfeab;
data_inb = 16'h49a;
#10;
address_ina = 198;
address_inb = 199;
data_ina = 16'h129;
data_inb = 16'hfa9b;
#10;
address_ina = 200;
address_inb = 201;
data_ina = 16'h1a8;
data_inb = 16'hfbed;
#10;
address_ina = 202;
address_inb = 203;
data_ina = 16'hfe31;
data_inb = 16'hfd60;
#10;
address_ina = 204;
address_inb = 205;
data_ina = 16'h333;
data_inb = 16'h538;
#10;
address_ina = 206;
address_inb = 207;
data_ina = 16'hfa45;
data_inb = 16'hfb91;
#10;
address_ina = 208;
address_inb = 209;
data_ina = 16'hff62;
data_inb = 16'hfbfe;
#10;
address_ina = 210;
address_inb = 211;
data_ina = 16'h344;
data_inb = 16'hfef2;
#10;
address_ina = 212;
address_inb = 213;
data_ina = 16'h61b;
data_inb = 16'hfec2;
#10;
address_ina = 214;
address_inb = 215;
data_ina = 16'hff97;
data_inb = 16'hfd80;
#10;
address_ina = 216;
address_inb = 217;
data_ina = 16'hff10;
data_inb = 16'hfb87;
#10;
address_ina = 218;
address_inb = 219;
data_ina = 16'hff3f;
data_inb = 16'h3e8;
#10;
address_ina = 220;
address_inb = 221;
data_ina = 16'hfdd9;
data_inb = 16'hfeec;
#10;
address_ina = 222;
address_inb = 223;
data_ina = 16'hfcf7;
data_inb = 16'hffbf;
#10;
address_ina = 224;
address_inb = 225;
data_ina = 16'hfc79;
data_inb = 16'h10c;
#10;
address_ina = 226;
address_inb = 227;
data_ina = 16'h5d1;
data_inb = 16'h26b;
#10;
address_ina = 228;
address_inb = 229;
data_ina = 16'h3be;
data_inb = 16'h4cb;
#10;
address_ina = 230;
address_inb = 231;
data_ina = 16'h119;
data_inb = 16'h436;
#10;
address_ina = 232;
address_inb = 233;
data_ina = 16'hfb68;
data_inb = 16'h4f8;
#10;
address_ina = 234;
address_inb = 235;
data_ina = 16'hfbf0;
data_inb = 16'h531;
#10;
address_ina = 236;
address_inb = 237;
data_ina = 16'hfd60;
data_inb = 16'hfccb;
#10;
address_ina = 238;
address_inb = 239;
data_ina = 16'h182;
data_inb = 16'h653;
#10;
address_ina = 240;
address_inb = 241;
data_ina = 16'hfe06;
data_inb = 16'hfe8b;
#10;
address_ina = 242;
address_inb = 243;
data_ina = 16'h393;
data_inb = 16'hfdaf;
#10;
address_ina = 244;
address_inb = 245;
data_ina = 16'hff9a;
data_inb = 16'hff80;
#10;
address_ina = 246;
address_inb = 247;
data_ina = 16'hfe05;
data_inb = 16'h133;
#10;
address_ina = 248;
address_inb = 249;
data_ina = 16'h323;
data_inb = 16'hfb1f;
#10;
address_ina = 250;
address_inb = 251;
data_ina = 16'hf9e8;
data_inb = 16'h2f7;
#10;
address_ina = 252;
address_inb = 253;
data_ina = 16'hfab4;
data_inb = 16'h39e;
#10;
address_ina = 254;
address_inb = 255;
data_ina = 16'hfeb3;
data_inb = 16'h268;
#10;
        wait(init_done);
        #30
        we = 0;
        // Start processing
         
		  #38000

        start = 0;



//        wait (wr_req);
//		  wait (!wr_req);
//		   rd_req = 1;
		  wait(done);
		  #20000
rd_req = 1;
        #70 
		  start = 1;
		 #80 
wait(rd_empty)
rd_req = 0;

$display("Finished the NTT test Number %d",test_num);
////Begin test number #59//////////////
rst = 1;

//#1000
start = 1;
mode = 1; //NTT 0 // INTT 1

// Reset for a few clock cycles

#1000

rst = 0;
test_num = test_num + 1;
#1000
we = 1;
address_ina = 0;
address_inb = 1;
data_ina = 16'hff7d;
data_inb = 16'h2c8;
#10;
address_ina = 2;
address_inb = 3;
data_ina = 16'hfcf9;
data_inb = 16'hfaa6;
#10;
address_ina = 4;
address_inb = 5;
data_ina = 16'h58;
data_inb = 16'h43c;
#10;
address_ina = 6;
address_inb = 7;
data_ina = 16'h23e;
data_inb = 16'hfaa2;
#10;
address_ina = 8;
address_inb = 9;
data_ina = 16'hff48;
data_inb = 16'h1dc;
#10;
address_ina = 10;
address_inb = 11;
data_ina = 16'h5d3;
data_inb = 16'hfdc0;
#10;
address_ina = 12;
address_inb = 13;
data_ina = 16'hfce1;
data_inb = 16'h5e1;
#10;
address_ina = 14;
address_inb = 15;
data_ina = 16'h66e;
data_inb = 16'h3c3;
#10;
address_ina = 16;
address_inb = 17;
data_ina = 16'hfe10;
data_inb = 16'hfb44;
#10;
address_ina = 18;
address_inb = 19;
data_ina = 16'h278;
data_inb = 16'hfbac;
#10;
address_ina = 20;
address_inb = 21;
data_ina = 16'hfe40;
data_inb = 16'h442;
#10;
address_ina = 22;
address_inb = 23;
data_ina = 16'hff62;
data_inb = 16'hfda7;
#10;
address_ina = 24;
address_inb = 25;
data_ina = 16'h4e;
data_inb = 16'heb;
#10;
address_ina = 26;
address_inb = 27;
data_ina = 16'h35e;
data_inb = 16'h26e;
#10;
address_ina = 28;
address_inb = 29;
data_ina = 16'hfc2c;
data_inb = 16'h4bb;
#10;
address_ina = 30;
address_inb = 31;
data_ina = 16'h28;
data_inb = 16'hfb60;
#10;
address_ina = 32;
address_inb = 33;
data_ina = 16'hfb1d;
data_inb = 16'h41d;
#10;
address_ina = 34;
address_inb = 35;
data_ina = 16'hfc79;
data_inb = 16'h426;
#10;
address_ina = 36;
address_inb = 37;
data_ina = 16'hfb75;
data_inb = 16'h193;
#10;
address_ina = 38;
address_inb = 39;
data_ina = 16'hfcc1;
data_inb = 16'hfeb0;
#10;
address_ina = 40;
address_inb = 41;
data_ina = 16'h164;
data_inb = 16'h5fa;
#10;
address_ina = 42;
address_inb = 43;
data_ina = 16'h37;
data_inb = 16'hfd86;
#10;
address_ina = 44;
address_inb = 45;
data_ina = 16'hfe9e;
data_inb = 16'hfee9;
#10;
address_ina = 46;
address_inb = 47;
data_ina = 16'h3f1;
data_inb = 16'h623;
#10;
address_ina = 48;
address_inb = 49;
data_ina = 16'hfd3e;
data_inb = 16'hfde8;
#10;
address_ina = 50;
address_inb = 51;
data_ina = 16'hfc89;
data_inb = 16'h4d8;
#10;
address_ina = 52;
address_inb = 53;
data_ina = 16'hfcbd;
data_inb = 16'hfb3b;
#10;
address_ina = 54;
address_inb = 55;
data_ina = 16'h609;
data_inb = 16'hfd3d;
#10;
address_ina = 56;
address_inb = 57;
data_ina = 16'h134;
data_inb = 16'hffe9;
#10;
address_ina = 58;
address_inb = 59;
data_ina = 16'hff64;
data_inb = 16'h29f;
#10;
address_ina = 60;
address_inb = 61;
data_ina = 16'h1ec;
data_inb = 16'h5c5;
#10;
address_ina = 62;
address_inb = 63;
data_ina = 16'h4fd;
data_inb = 16'h187;
#10;
address_ina = 64;
address_inb = 65;
data_ina = 16'hf9e4;
data_inb = 16'h303;
#10;
address_ina = 66;
address_inb = 67;
data_ina = 16'h40f;
data_inb = 16'h13d;
#10;
address_ina = 68;
address_inb = 69;
data_ina = 16'hff29;
data_inb = 16'h2c9;
#10;
address_ina = 70;
address_inb = 71;
data_ina = 16'hfec9;
data_inb = 16'hfec0;
#10;
address_ina = 72;
address_inb = 73;
data_ina = 16'hfde5;
data_inb = 16'hfdaa;
#10;
address_ina = 74;
address_inb = 75;
data_ina = 16'h258;
data_inb = 16'hfc14;
#10;
address_ina = 76;
address_inb = 77;
data_ina = 16'h434;
data_inb = 16'hf9f7;
#10;
address_ina = 78;
address_inb = 79;
data_ina = 16'hff65;
data_inb = 16'hff04;
#10;
address_ina = 80;
address_inb = 81;
data_ina = 16'hfdcb;
data_inb = 16'hf9b4;
#10;
address_ina = 82;
address_inb = 83;
data_ina = 16'h163;
data_inb = 16'hfcf2;
#10;
address_ina = 84;
address_inb = 85;
data_ina = 16'h602;
data_inb = 16'hfd73;
#10;
address_ina = 86;
address_inb = 87;
data_ina = 16'hfa17;
data_inb = 16'h384;
#10;
address_ina = 88;
address_inb = 89;
data_ina = 16'h2c6;
data_inb = 16'h323;
#10;
address_ina = 90;
address_inb = 91;
data_ina = 16'h3d;
data_inb = 16'hfeb5;
#10;
address_ina = 92;
address_inb = 93;
data_ina = 16'h331;
data_inb = 16'h367;
#10;
address_ina = 94;
address_inb = 95;
data_ina = 16'hfaa2;
data_inb = 16'hfcd6;
#10;
address_ina = 96;
address_inb = 97;
data_ina = 16'hfad8;
data_inb = 16'h3b2;
#10;
address_ina = 98;
address_inb = 99;
data_ina = 16'h1a9;
data_inb = 16'h568;
#10;
address_ina = 100;
address_inb = 101;
data_ina = 16'hfdb5;
data_inb = 16'hfa87;
#10;
address_ina = 102;
address_inb = 103;
data_ina = 16'h46;
data_inb = 16'hfc3a;
#10;
address_ina = 104;
address_inb = 105;
data_ina = 16'h1ec;
data_inb = 16'h18a;
#10;
address_ina = 106;
address_inb = 107;
data_ina = 16'h436;
data_inb = 16'hf9b2;
#10;
address_ina = 108;
address_inb = 109;
data_ina = 16'hff99;
data_inb = 16'h2d2;
#10;
address_ina = 110;
address_inb = 111;
data_ina = 16'hffee;
data_inb = 16'h30f;
#10;
address_ina = 112;
address_inb = 113;
data_ina = 16'h1f1;
data_inb = 16'hfda7;
#10;
address_ina = 114;
address_inb = 115;
data_ina = 16'h609;
data_inb = 16'h4f9;
#10;
address_ina = 116;
address_inb = 117;
data_ina = 16'hfa84;
data_inb = 16'hff22;
#10;
address_ina = 118;
address_inb = 119;
data_ina = 16'hfd67;
data_inb = 16'h319;
#10;
address_ina = 120;
address_inb = 121;
data_ina = 16'hfb17;
data_inb = 16'hfa43;
#10;
address_ina = 122;
address_inb = 123;
data_ina = 16'h4e0;
data_inb = 16'h2e7;
#10;
address_ina = 124;
address_inb = 125;
data_ina = 16'hfb5d;
data_inb = 16'hfe49;
#10;
address_ina = 126;
address_inb = 127;
data_ina = 16'h384;
data_inb = 16'h395;
#10;
address_ina = 128;
address_inb = 129;
data_ina = 16'h160;
data_inb = 16'hffff;
#10;
address_ina = 130;
address_inb = 131;
data_ina = 16'h390;
data_inb = 16'h2f1;
#10;
address_ina = 132;
address_inb = 133;
data_ina = 16'h4aa;
data_inb = 16'hf9c6;
#10;
address_ina = 134;
address_inb = 135;
data_ina = 16'hfe46;
data_inb = 16'hfefb;
#10;
address_ina = 136;
address_inb = 137;
data_ina = 16'hfd0e;
data_inb = 16'h217;
#10;
address_ina = 138;
address_inb = 139;
data_ina = 16'hfc8f;
data_inb = 16'h321;
#10;
address_ina = 140;
address_inb = 141;
data_ina = 16'h467;
data_inb = 16'hfd70;
#10;
address_ina = 142;
address_inb = 143;
data_ina = 16'h1db;
data_inb = 16'h628;
#10;
address_ina = 144;
address_inb = 145;
data_ina = 16'h5ba;
data_inb = 16'h421;
#10;
address_ina = 146;
address_inb = 147;
data_ina = 16'hfc1f;
data_inb = 16'hffeb;
#10;
address_ina = 148;
address_inb = 149;
data_ina = 16'hfd0e;
data_inb = 16'h455;
#10;
address_ina = 150;
address_inb = 151;
data_ina = 16'hfa41;
data_inb = 16'h182;
#10;
address_ina = 152;
address_inb = 153;
data_ina = 16'hfd94;
data_inb = 16'hfc0f;
#10;
address_ina = 154;
address_inb = 155;
data_ina = 16'hfe8e;
data_inb = 16'hfb66;
#10;
address_ina = 156;
address_inb = 157;
data_ina = 16'h4d7;
data_inb = 16'h27f;
#10;
address_ina = 158;
address_inb = 159;
data_ina = 16'h17f;
data_inb = 16'hab;
#10;
address_ina = 160;
address_inb = 161;
data_ina = 16'h36a;
data_inb = 16'hea;
#10;
address_ina = 162;
address_inb = 163;
data_ina = 16'ha1;
data_inb = 16'h467;
#10;
address_ina = 164;
address_inb = 165;
data_ina = 16'h2ed;
data_inb = 16'h53a;
#10;
address_ina = 166;
address_inb = 167;
data_ina = 16'h68;
data_inb = 16'hfc9c;
#10;
address_ina = 168;
address_inb = 169;
data_ina = 16'hfc4d;
data_inb = 16'h578;
#10;
address_ina = 170;
address_inb = 171;
data_ina = 16'h34f;
data_inb = 16'h5a4;
#10;
address_ina = 172;
address_inb = 173;
data_ina = 16'hab;
data_inb = 16'hfc2e;
#10;
address_ina = 174;
address_inb = 175;
data_ina = 16'hfc13;
data_inb = 16'hfec2;
#10;
address_ina = 176;
address_inb = 177;
data_ina = 16'h1af;
data_inb = 16'hfa73;
#10;
address_ina = 178;
address_inb = 179;
data_ina = 16'hfc44;
data_inb = 16'hfb6c;
#10;
address_ina = 180;
address_inb = 181;
data_ina = 16'h541;
data_inb = 16'hfe84;
#10;
address_ina = 182;
address_inb = 183;
data_ina = 16'h359;
data_inb = 16'h24c;
#10;
address_ina = 184;
address_inb = 185;
data_ina = 16'hfe2b;
data_inb = 16'h2b;
#10;
address_ina = 186;
address_inb = 187;
data_ina = 16'hfcf9;
data_inb = 16'h4f5;
#10;
address_ina = 188;
address_inb = 189;
data_ina = 16'h66d;
data_inb = 16'hff69;
#10;
address_ina = 190;
address_inb = 191;
data_ina = 16'hfd47;
data_inb = 16'h3f;
#10;
address_ina = 192;
address_inb = 193;
data_ina = 16'h18a;
data_inb = 16'hfa8d;
#10;
address_ina = 194;
address_inb = 195;
data_ina = 16'h4cd;
data_inb = 16'hf9;
#10;
address_ina = 196;
address_inb = 197;
data_ina = 16'h331;
data_inb = 16'hfb91;
#10;
address_ina = 198;
address_inb = 199;
data_ina = 16'h38a;
data_inb = 16'h362;
#10;
address_ina = 200;
address_inb = 201;
data_ina = 16'h18d;
data_inb = 16'h680;
#10;
address_ina = 202;
address_inb = 203;
data_ina = 16'hfb3f;
data_inb = 16'hfb64;
#10;
address_ina = 204;
address_inb = 205;
data_ina = 16'hfe83;
data_inb = 16'h42b;
#10;
address_ina = 206;
address_inb = 207;
data_ina = 16'hfa1b;
data_inb = 16'h59c;
#10;
address_ina = 208;
address_inb = 209;
data_ina = 16'hffe5;
data_inb = 16'h586;
#10;
address_ina = 210;
address_inb = 211;
data_ina = 16'h374;
data_inb = 16'hd6;
#10;
address_ina = 212;
address_inb = 213;
data_ina = 16'h74;
data_inb = 16'hfba6;
#10;
address_ina = 214;
address_inb = 215;
data_ina = 16'h4c3;
data_inb = 16'h34f;
#10;
address_ina = 216;
address_inb = 217;
data_ina = 16'h41c;
data_inb = 16'h2f;
#10;
address_ina = 218;
address_inb = 219;
data_ina = 16'h27e;
data_inb = 16'h3b5;
#10;
address_ina = 220;
address_inb = 221;
data_ina = 16'hff7e;
data_inb = 16'h61d;
#10;
address_ina = 222;
address_inb = 223;
data_ina = 16'hfd37;
data_inb = 16'hfed3;
#10;
address_ina = 224;
address_inb = 225;
data_ina = 16'h2fe;
data_inb = 16'hfb53;
#10;
address_ina = 226;
address_inb = 227;
data_ina = 16'hfe14;
data_inb = 16'hfb9c;
#10;
address_ina = 228;
address_inb = 229;
data_ina = 16'hfdeb;
data_inb = 16'h347;
#10;
address_ina = 230;
address_inb = 231;
data_ina = 16'hfcf9;
data_inb = 16'h575;
#10;
address_ina = 232;
address_inb = 233;
data_ina = 16'h549;
data_inb = 16'h163;
#10;
address_ina = 234;
address_inb = 235;
data_ina = 16'hfd8c;
data_inb = 16'hfae2;
#10;
address_ina = 236;
address_inb = 237;
data_ina = 16'h5cc;
data_inb = 16'h2e;
#10;
address_ina = 238;
address_inb = 239;
data_ina = 16'h397;
data_inb = 16'hfab9;
#10;
address_ina = 240;
address_inb = 241;
data_ina = 16'h1bb;
data_inb = 16'h24;
#10;
address_ina = 242;
address_inb = 243;
data_ina = 16'hff1d;
data_inb = 16'hf9a0;
#10;
address_ina = 244;
address_inb = 245;
data_ina = 16'h651;
data_inb = 16'hfb13;
#10;
address_ina = 246;
address_inb = 247;
data_ina = 16'h5f8;
data_inb = 16'hfb03;
#10;
address_ina = 248;
address_inb = 249;
data_ina = 16'hfd74;
data_inb = 16'h142;
#10;
address_ina = 250;
address_inb = 251;
data_ina = 16'h566;
data_inb = 16'hfa6a;
#10;
address_ina = 252;
address_inb = 253;
data_ina = 16'hff97;
data_inb = 16'hfd24;
#10;
address_ina = 254;
address_inb = 255;
data_ina = 16'h2a0;
data_inb = 16'h5ef;
#10;
        wait(init_done);
        #30
        we = 0;
        // Start processing
         
		  #38000

        start = 0;



//        wait (wr_req);
//		  wait (!wr_req);
//		   rd_req = 1;
		  wait(done);
		  #20000
rd_req = 1;
        #70 
		  start = 1;
		 #80 
wait(rd_empty)
rd_req = 0;

$display("Finished the NTT test Number %d",test_num);
////Begin test number #60//////////////
rst = 1;

//#1000
start = 1;
mode = 0; //NTT 0 // INTT 1

// Reset for a few clock cycles

#1000

rst = 0;
test_num = test_num + 1;
#1000
we = 1;
address_ina = 0;
address_inb = 1;
data_ina = 16'h656;
data_inb = 16'hb19;
#10;
address_ina = 2;
address_inb = 3;
data_ina = 16'h166;
data_inb = 16'h1f1;
#10;
address_ina = 4;
address_inb = 5;
data_ina = 16'hbb9;
data_inb = 16'h851;
#10;
address_ina = 6;
address_inb = 7;
data_ina = 16'hb9f;
data_inb = 16'h6c8;
#10;
address_ina = 8;
address_inb = 9;
data_ina = 16'h38b;
data_inb = 16'h23f;
#10;
address_ina = 10;
address_inb = 11;
data_ina = 16'h3c9;
data_inb = 16'ha08;
#10;
address_ina = 12;
address_inb = 13;
data_ina = 16'h6e5;
data_inb = 16'h559;
#10;
address_ina = 14;
address_inb = 15;
data_ina = 16'h84e;
data_inb = 16'h3b5;
#10;
address_ina = 16;
address_inb = 17;
data_ina = 16'h5fb;
data_inb = 16'h92e;
#10;
address_ina = 18;
address_inb = 19;
data_ina = 16'h3f3;
data_inb = 16'h45b;
#10;
address_ina = 20;
address_inb = 21;
data_ina = 16'h2c1;
data_inb = 16'h7c;
#10;
address_ina = 22;
address_inb = 23;
data_ina = 16'h586;
data_inb = 16'h767;
#10;
address_ina = 24;
address_inb = 25;
data_ina = 16'haa1;
data_inb = 16'ha74;
#10;
address_ina = 26;
address_inb = 27;
data_ina = 16'ha67;
data_inb = 16'hb2a;
#10;
address_ina = 28;
address_inb = 29;
data_ina = 16'h36e;
data_inb = 16'h193;
#10;
address_ina = 30;
address_inb = 31;
data_ina = 16'hbbf;
data_inb = 16'h159;
#10;
address_ina = 32;
address_inb = 33;
data_ina = 16'h1e8;
data_inb = 16'hf1;
#10;
address_ina = 34;
address_inb = 35;
data_ina = 16'h52e;
data_inb = 16'hcd;
#10;
address_ina = 36;
address_inb = 37;
data_ina = 16'h9d8;
data_inb = 16'h5ee;
#10;
address_ina = 38;
address_inb = 39;
data_ina = 16'h49f;
data_inb = 16'h4d0;
#10;
address_ina = 40;
address_inb = 41;
data_ina = 16'h865;
data_inb = 16'hb3d;
#10;
address_ina = 42;
address_inb = 43;
data_ina = 16'h3ed;
data_inb = 16'h35e;
#10;
address_ina = 44;
address_inb = 45;
data_ina = 16'ha94;
data_inb = 16'h44e;
#10;
address_ina = 46;
address_inb = 47;
data_ina = 16'h986;
data_inb = 16'h6b8;
#10;
address_ina = 48;
address_inb = 49;
data_ina = 16'hae2;
data_inb = 16'h19d;
#10;
address_ina = 50;
address_inb = 51;
data_ina = 16'h19d;
data_inb = 16'h89c;
#10;
address_ina = 52;
address_inb = 53;
data_ina = 16'ha9b;
data_inb = 16'h2ab;
#10;
address_ina = 54;
address_inb = 55;
data_ina = 16'hbfa;
data_inb = 16'h8f1;
#10;
address_ina = 56;
address_inb = 57;
data_ina = 16'h44e;
data_inb = 16'h47c;
#10;
address_ina = 58;
address_inb = 59;
data_ina = 16'h4ca;
data_inb = 16'hac5;
#10;
address_ina = 60;
address_inb = 61;
data_ina = 16'h344;
data_inb = 16'h246;
#10;
address_ina = 62;
address_inb = 63;
data_ina = 16'h726;
data_inb = 16'h62;
#10;
address_ina = 64;
address_inb = 65;
data_ina = 16'h68;
data_inb = 16'h74d;
#10;
address_ina = 66;
address_inb = 67;
data_ina = 16'h5f5;
data_inb = 16'hafc;
#10;
address_ina = 68;
address_inb = 69;
data_ina = 16'h5ad;
data_inb = 16'hce4;
#10;
address_ina = 70;
address_inb = 71;
data_ina = 16'h179;
data_inb = 16'h17;
#10;
address_ina = 72;
address_inb = 73;
data_ina = 16'h8f1;
data_inb = 16'hc03;
#10;
address_ina = 74;
address_inb = 75;
data_ina = 16'hb16;
data_inb = 16'hc4e;
#10;
address_ina = 76;
address_inb = 77;
data_ina = 16'hbbc;
data_inb = 16'h26d;
#10;
address_ina = 78;
address_inb = 79;
data_ina = 16'h697;
data_inb = 16'h31;
#10;
address_ina = 80;
address_inb = 81;
data_ina = 16'ha08;
data_inb = 16'h67d;
#10;
address_ina = 82;
address_inb = 83;
data_ina = 16'h528;
data_inb = 16'h79f;
#10;
address_ina = 84;
address_inb = 85;
data_ina = 16'hc31;
data_inb = 16'hc44;
#10;
address_ina = 86;
address_inb = 87;
data_ina = 16'h496;
data_inb = 16'h6ec;
#10;
address_ina = 88;
address_inb = 89;
data_ina = 16'h81d;
data_inb = 16'h5a7;
#10;
address_ina = 90;
address_inb = 91;
data_ina = 16'h249;
data_inb = 16'hc58;
#10;
address_ina = 92;
address_inb = 93;
data_ina = 16'h2b8;
data_inb = 16'h1d;
#10;
address_ina = 94;
address_inb = 95;
data_ina = 16'hc5b;
data_inb = 16'hbd3;
#10;
address_ina = 96;
address_inb = 97;
data_ina = 16'h892;
data_inb = 16'hb03;
#10;
address_ina = 98;
address_inb = 99;
data_ina = 16'h6be;
data_inb = 16'h222;
#10;
address_ina = 100;
address_inb = 101;
data_ina = 16'hb6;
data_inb = 16'h726;
#10;
address_ina = 102;
address_inb = 103;
data_ina = 16'hb61;
data_inb = 16'h79f;
#10;
address_ina = 104;
address_inb = 105;
data_ina = 16'h48;
data_inb = 16'h8c;
#10;
address_ina = 106;
address_inb = 107;
data_ina = 16'hbe9;
data_inb = 16'h294;
#10;
address_ina = 108;
address_inb = 109;
data_ina = 16'h81d;
data_inb = 16'h448;
#10;
address_ina = 110;
address_inb = 111;
data_ina = 16'h803;
data_inb = 16'ha02;
#10;
address_ina = 112;
address_inb = 113;
data_ina = 16'h8f1;
data_inb = 16'h3b;
#10;
address_ina = 114;
address_inb = 115;
data_ina = 16'h1b7;
data_inb = 16'h3ac;
#10;
address_ina = 116;
address_inb = 117;
data_ina = 16'h90e;
data_inb = 16'h85;
#10;
address_ina = 118;
address_inb = 119;
data_ina = 16'hc9c;
data_inb = 16'h3ed;
#10;
address_ina = 120;
address_inb = 121;
data_ina = 16'h7b2;
data_inb = 16'hab5;
#10;
address_ina = 122;
address_inb = 123;
data_ina = 16'h1ce;
data_inb = 16'h6d2;
#10;
address_ina = 124;
address_inb = 125;
data_ina = 16'h8ed;
data_inb = 16'hb81;
#10;
address_ina = 126;
address_inb = 127;
data_ina = 16'h5b4;
data_inb = 16'h270;
#10;
address_ina = 128;
address_inb = 129;
data_ina = 16'h444;
data_inb = 16'h821;
#10;
address_ina = 130;
address_inb = 131;
data_ina = 16'hb23;
data_inb = 16'h990;
#10;
address_ina = 132;
address_inb = 133;
data_ina = 16'h555;
data_inb = 16'ha60;
#10;
address_ina = 134;
address_inb = 135;
data_ina = 16'ha87;
data_inb = 16'h44;
#10;
address_ina = 136;
address_inb = 137;
data_ina = 16'h347;
data_inb = 16'h58;
#10;
address_ina = 138;
address_inb = 139;
data_ina = 16'h781;
data_inb = 16'ha7a;
#10;
address_ina = 140;
address_inb = 141;
data_ina = 16'h41a;
data_inb = 16'h952;
#10;
address_ina = 142;
address_inb = 143;
data_ina = 16'h41;
data_inb = 16'h5b0;
#10;
address_ina = 144;
address_inb = 145;
data_ina = 16'hcda;
data_inb = 16'hb33;
#10;
address_ina = 146;
address_inb = 147;
data_ina = 16'h455;
data_inb = 16'h7c2;
#10;
address_ina = 148;
address_inb = 149;
data_ina = 16'h84b;
data_inb = 16'h33d;
#10;
address_ina = 150;
address_inb = 151;
data_ina = 16'h15c;
data_inb = 16'ha3;
#10;
address_ina = 152;
address_inb = 153;
data_ina = 16'h6e9;
data_inb = 16'h542;
#10;
address_ina = 154;
address_inb = 155;
data_ina = 16'hb23;
data_inb = 16'h212;
#10;
address_ina = 156;
address_inb = 157;
data_ina = 16'h385;
data_inb = 16'h2e2;
#10;
address_ina = 158;
address_inb = 159;
data_ina = 16'hc27;
data_inb = 16'h414;
#10;
address_ina = 160;
address_inb = 161;
data_ina = 16'h593;
data_inb = 16'h84e;
#10;
address_ina = 162;
address_inb = 163;
data_ina = 16'haf6;
data_inb = 16'h2d5;
#10;
address_ina = 164;
address_inb = 165;
data_ina = 16'h709;
data_inb = 16'h4bd;
#10;
address_ina = 166;
address_inb = 167;
data_ina = 16'haef;
data_inb = 16'h1e8;
#10;
address_ina = 168;
address_inb = 169;
data_ina = 16'ha39;
data_inb = 16'h36e;
#10;
address_ina = 170;
address_inb = 171;
data_ina = 16'h4a3;
data_inb = 16'h326;
#10;
address_ina = 172;
address_inb = 173;
data_ina = 16'hce4;
data_inb = 16'h478;
#10;
address_ina = 174;
address_inb = 175;
data_ina = 16'h82;
data_inb = 16'h589;
#10;
address_ina = 176;
address_inb = 177;
data_ina = 16'h492;
data_inb = 16'h155;
#10;
address_ina = 178;
address_inb = 179;
data_ina = 16'h52b;
data_inb = 16'h6d8;
#10;
address_ina = 180;
address_inb = 181;
data_ina = 16'h5b7;
data_inb = 16'hc27;
#10;
address_ina = 182;
address_inb = 183;
data_ina = 16'h1ee;
data_inb = 16'hca;
#10;
address_ina = 184;
address_inb = 185;
data_ina = 16'h7ac;
data_inb = 16'h38b;
#10;
address_ina = 186;
address_inb = 187;
data_ina = 16'h778;
data_inb = 16'hca3;
#10;
address_ina = 188;
address_inb = 189;
data_ina = 16'hae9;
data_inb = 16'hc41;
#10;
address_ina = 190;
address_inb = 191;
data_ina = 16'h618;
data_inb = 16'ha81;
#10;
address_ina = 192;
address_inb = 193;
data_ina = 16'h8e0;
data_inb = 16'hb3d;
#10;
address_ina = 194;
address_inb = 195;
data_ina = 16'h2d8;
data_inb = 16'h9c4;
#10;
address_ina = 196;
address_inb = 197;
data_ina = 16'ha8a;
data_inb = 16'h710;
#10;
address_ina = 198;
address_inb = 199;
data_ina = 16'h851;
data_inb = 16'h186;
#10;
address_ina = 200;
address_inb = 201;
data_ina = 16'h3cf;
data_inb = 16'h1c7;
#10;
address_ina = 202;
address_inb = 203;
data_ina = 16'h798;
data_inb = 16'h2c5;
#10;
address_ina = 204;
address_inb = 205;
data_ina = 16'h77e;
data_inb = 16'hb26;
#10;
address_ina = 206;
address_inb = 207;
data_ina = 16'h34d;
data_inb = 16'h414;
#10;
address_ina = 208;
address_inb = 209;
data_ina = 16'hafc;
data_inb = 16'h5b;
#10;
address_ina = 210;
address_inb = 211;
data_ina = 16'h5ca;
data_inb = 16'hc3b;
#10;
address_ina = 212;
address_inb = 213;
data_ina = 16'h72;
data_inb = 16'hbcc;
#10;
address_ina = 214;
address_inb = 215;
data_ina = 16'hcdd;
data_inb = 16'h12b;
#10;
address_ina = 216;
address_inb = 217;
data_ina = 16'h618;
data_inb = 16'h424;
#10;
address_ina = 218;
address_inb = 219;
data_ina = 16'h56c;
data_inb = 16'h1aa;
#10;
address_ina = 220;
address_inb = 221;
data_ina = 16'h249;
data_inb = 16'h3bf;
#10;
address_ina = 222;
address_inb = 223;
data_ina = 16'h81d;
data_inb = 16'hd7;
#10;
address_ina = 224;
address_inb = 225;
data_ina = 16'hcd3;
data_inb = 16'ha53;
#10;
address_ina = 226;
address_inb = 227;
data_ina = 16'h364;
data_inb = 16'h48f;
#10;
address_ina = 228;
address_inb = 229;
data_ina = 16'hbb5;
data_inb = 16'h6d2;
#10;
address_ina = 230;
address_inb = 231;
data_ina = 16'h138;
data_inb = 16'h414;
#10;
address_ina = 232;
address_inb = 233;
data_ina = 16'h294;
data_inb = 16'h6c2;
#10;
address_ina = 234;
address_inb = 235;
data_ina = 16'h643;
data_inb = 16'h67d;
#10;
address_ina = 236;
address_inb = 237;
data_ina = 16'h388;
data_inb = 16'hadf;
#10;
address_ina = 238;
address_inb = 239;
data_ina = 16'h663;
data_inb = 16'h371;
#10;
address_ina = 240;
address_inb = 241;
data_ina = 16'h58;
data_inb = 16'h62;
#10;
address_ina = 242;
address_inb = 243;
data_ina = 16'h53b;
data_inb = 16'h810;
#10;
address_ina = 244;
address_inb = 245;
data_ina = 16'h817;
data_inb = 16'hccd;
#10;
address_ina = 246;
address_inb = 247;
data_ina = 16'h2f2;
data_inb = 16'h61c;
#10;
address_ina = 248;
address_inb = 249;
data_ina = 16'h4ea;
data_inb = 16'ha74;
#10;
address_ina = 250;
address_inb = 251;
data_ina = 16'h892;
data_inb = 16'h138;
#10;
address_ina = 252;
address_inb = 253;
data_ina = 16'h656;
data_inb = 16'h47c;
#10;
address_ina = 254;
address_inb = 255;
data_ina = 16'h7a5;
data_inb = 16'h86f;
#10;
        wait(init_done);
        #30
        we = 0;
        // Start processing
         
		  #38000

        start = 0;



//        wait (wr_req);
//		  wait (!wr_req);
//		   rd_req = 1;
		  wait(done);
		  #20000
rd_req = 1;
        #70 
		  start = 1;
		 #80 
wait(rd_empty)
rd_req = 0;

$display("Finished the NTT test Number %d",test_num);
////Begin test number #61//////////////
rst = 1;

//#1000
start = 1;
mode = 0; //NTT 0 // INTT 1

// Reset for a few clock cycles

#1000

rst = 0;
test_num = test_num + 1;
#1000
we = 1;
address_ina = 0;
address_inb = 1;
data_ina = 16'h414;
data_inb = 16'h6d5;
#10;
address_ina = 2;
address_inb = 3;
data_ina = 16'h959;
data_inb = 16'h52e;
#10;
address_ina = 4;
address_inb = 5;
data_ina = 16'h562;
data_inb = 16'h5f5;
#10;
address_ina = 6;
address_inb = 7;
data_ina = 16'h5f8;
data_inb = 16'hcfa;
#10;
address_ina = 8;
address_inb = 9;
data_ina = 16'h79f;
data_inb = 16'h5ba;
#10;
address_ina = 10;
address_inb = 11;
data_ina = 16'h656;
data_inb = 16'h169;
#10;
address_ina = 12;
address_inb = 13;
data_ina = 16'h7b9;
data_inb = 16'h79b;
#10;
address_ina = 14;
address_inb = 15;
data_ina = 16'h306;
data_inb = 16'h6d5;
#10;
address_ina = 16;
address_inb = 17;
data_ina = 16'hbe3;
data_inb = 16'h111;
#10;
address_ina = 18;
address_inb = 19;
data_ina = 16'h744;
data_inb = 16'h45e;
#10;
address_ina = 20;
address_inb = 21;
data_ina = 16'hb67;
data_inb = 16'h78e;
#10;
address_ina = 22;
address_inb = 23;
data_ina = 16'h6be;
data_inb = 16'hc37;
#10;
address_ina = 24;
address_inb = 25;
data_ina = 16'hb9b;
data_inb = 16'h26d;
#10;
address_ina = 26;
address_inb = 27;
data_ina = 16'h88c;
data_inb = 16'hc2a;
#10;
address_ina = 28;
address_inb = 29;
data_ina = 16'hcbd;
data_inb = 16'h521;
#10;
address_ina = 30;
address_inb = 31;
data_ina = 16'ha1c;
data_inb = 16'h3c2;
#10;
address_ina = 32;
address_inb = 33;
data_ina = 16'h424;
data_inb = 16'h2c8;
#10;
address_ina = 34;
address_inb = 35;
data_ina = 16'h319;
data_inb = 16'h2d5;
#10;
address_ina = 36;
address_inb = 37;
data_ina = 16'h737;
data_inb = 16'h4a3;
#10;
address_ina = 38;
address_inb = 39;
data_ina = 16'hb92;
data_inb = 16'h92;
#10;
address_ina = 40;
address_inb = 41;
data_ina = 16'hac2;
data_inb = 16'h7;
#10;
address_ina = 42;
address_inb = 43;
data_ina = 16'h287;
data_inb = 16'h465;
#10;
address_ina = 44;
address_inb = 45;
data_ina = 16'h6ff;
data_inb = 16'h9ff;
#10;
address_ina = 46;
address_inb = 47;
data_ina = 16'h5ca;
data_inb = 16'h69b;
#10;
address_ina = 48;
address_inb = 49;
data_ina = 16'h8c3;
data_inb = 16'h952;
#10;
address_ina = 50;
address_inb = 51;
data_ina = 16'hdd;
data_inb = 16'h660;
#10;
address_ina = 52;
address_inb = 53;
data_ina = 16'h9c7;
data_inb = 16'hac;
#10;
address_ina = 54;
address_inb = 55;
data_ina = 16'h1f8;
data_inb = 16'hb3a;
#10;
address_ina = 56;
address_inb = 57;
data_ina = 16'h579;
data_inb = 16'hbd3;
#10;
address_ina = 58;
address_inb = 59;
data_ina = 16'haa4;
data_inb = 16'h562;
#10;
address_ina = 60;
address_inb = 61;
data_ina = 16'h2ab;
data_inb = 16'h42e;
#10;
address_ina = 62;
address_inb = 63;
data_ina = 16'h96;
data_inb = 16'hdd;
#10;
address_ina = 64;
address_inb = 65;
data_ina = 16'h183;
data_inb = 16'h407;
#10;
address_ina = 66;
address_inb = 67;
data_ina = 16'h2c1;
data_inb = 16'h4e0;
#10;
address_ina = 68;
address_inb = 69;
data_ina = 16'h6cb;
data_inb = 16'h9e8;
#10;
address_ina = 70;
address_inb = 71;
data_ina = 16'h2c5;
data_inb = 16'h945;
#10;
address_ina = 72;
address_inb = 73;
data_ina = 16'h7;
data_inb = 16'hb26;
#10;
address_ina = 74;
address_inb = 75;
data_ina = 16'h354;
data_inb = 16'h788;
#10;
address_ina = 76;
address_inb = 77;
data_ina = 16'h80a;
data_inb = 16'h4b0;
#10;
address_ina = 78;
address_inb = 79;
data_ina = 16'h1f5;
data_inb = 16'h414;
#10;
address_ina = 80;
address_inb = 81;
data_ina = 16'hcc0;
data_inb = 16'h528;
#10;
address_ina = 82;
address_inb = 83;
data_ina = 16'h969;
data_inb = 16'h280;
#10;
address_ina = 84;
address_inb = 85;
data_ina = 16'h72;
data_inb = 16'hb88;
#10;
address_ina = 86;
address_inb = 87;
data_ina = 16'h878;
data_inb = 16'h3e6;
#10;
address_ina = 88;
address_inb = 89;
data_ina = 16'h901;
data_inb = 16'hcf7;
#10;
address_ina = 90;
address_inb = 91;
data_ina = 16'hba5;
data_inb = 16'h8f;
#10;
address_ina = 92;
address_inb = 93;
data_ina = 16'hccd;
data_inb = 16'hca6;
#10;
address_ina = 94;
address_inb = 95;
data_ina = 16'h1b7;
data_inb = 16'h5b0;
#10;
address_ina = 96;
address_inb = 97;
data_ina = 16'h2e2;
data_inb = 16'hb5e;
#10;
address_ina = 98;
address_inb = 99;
data_ina = 16'h4ed;
data_inb = 16'h629;
#10;
address_ina = 100;
address_inb = 101;
data_ina = 16'ha9;
data_inb = 16'h3fd;
#10;
address_ina = 102;
address_inb = 103;
data_ina = 16'h2a1;
data_inb = 16'hf1;
#10;
address_ina = 104;
address_inb = 105;
data_ina = 16'h904;
data_inb = 16'h8c0;
#10;
address_ina = 106;
address_inb = 107;
data_ina = 16'hb1d;
data_inb = 16'h716;
#10;
address_ina = 108;
address_inb = 109;
data_ina = 16'h45b;
data_inb = 16'h98d;
#10;
address_ina = 110;
address_inb = 111;
data_ina = 16'h650;
data_inb = 16'h73a;
#10;
address_ina = 112;
address_inb = 113;
data_ina = 16'h9ba;
data_inb = 16'h559;
#10;
address_ina = 114;
address_inb = 115;
data_ina = 16'h7c;
data_inb = 16'hba5;
#10;
address_ina = 116;
address_inb = 117;
data_ina = 16'h66a;
data_inb = 16'hc3;
#10;
address_ina = 118;
address_inb = 119;
data_ina = 16'h169;
data_inb = 16'h44b;
#10;
address_ina = 120;
address_inb = 121;
data_ina = 16'h55f;
data_inb = 16'h848;
#10;
address_ina = 122;
address_inb = 123;
data_ina = 16'h99;
data_inb = 16'h80d;
#10;
address_ina = 124;
address_inb = 125;
data_ina = 16'h22f;
data_inb = 16'h6a8;
#10;
address_ina = 126;
address_inb = 127;
data_ina = 16'hb57;
data_inb = 16'h7c2;
#10;
address_ina = 128;
address_inb = 129;
data_ina = 16'hc1a;
data_inb = 16'ha63;
#10;
address_ina = 130;
address_inb = 131;
data_ina = 16'h9c1;
data_inb = 16'hc3;
#10;
address_ina = 132;
address_inb = 133;
data_ina = 16'h21;
data_inb = 16'ha8a;
#10;
address_ina = 134;
address_inb = 135;
data_ina = 16'h3;
data_inb = 16'h37;
#10;
address_ina = 136;
address_inb = 137;
data_ina = 16'hea;
data_inb = 16'h9b0;
#10;
address_ina = 138;
address_inb = 139;
data_ina = 16'h785;
data_inb = 16'h94f;
#10;
address_ina = 140;
address_inb = 141;
data_ina = 16'h437;
data_inb = 16'h3af;
#10;
address_ina = 142;
address_inb = 143;
data_ina = 16'haff;
data_inb = 16'h9e1;
#10;
address_ina = 144;
address_inb = 145;
data_ina = 16'h75e;
data_inb = 16'hbf0;
#10;
address_ina = 146;
address_inb = 147;
data_ina = 16'h270;
data_inb = 16'h1d7;
#10;
address_ina = 148;
address_inb = 149;
data_ina = 16'h381;
data_inb = 16'h6d2;
#10;
address_ina = 150;
address_inb = 151;
data_ina = 16'h9db;
data_inb = 16'h57c;
#10;
address_ina = 152;
address_inb = 153;
data_ina = 16'h91e;
data_inb = 16'h518;
#10;
address_ina = 154;
address_inb = 155;
data_ina = 16'hb67;
data_inb = 16'h51;
#10;
address_ina = 156;
address_inb = 157;
data_ina = 16'ha6;
data_inb = 16'h29e;
#10;
address_ina = 158;
address_inb = 159;
data_ina = 16'hac2;
data_inb = 16'h625;
#10;
address_ina = 160;
address_inb = 161;
data_ina = 16'ha84;
data_inb = 16'h89c;
#10;
address_ina = 162;
address_inb = 163;
data_ina = 16'h12b;
data_inb = 16'hb6;
#10;
address_ina = 164;
address_inb = 165;
data_ina = 16'h6c8;
data_inb = 16'h10e;
#10;
address_ina = 166;
address_inb = 167;
data_ina = 16'hce4;
data_inb = 16'h53f;
#10;
address_ina = 168;
address_inb = 169;
data_ina = 16'h9d1;
data_inb = 16'hc7f;
#10;
address_ina = 170;
address_inb = 171;
data_ina = 16'h48c;
data_inb = 16'h993;
#10;
address_ina = 172;
address_inb = 173;
data_ina = 16'h80a;
data_inb = 16'haf9;
#10;
address_ina = 174;
address_inb = 175;
data_ina = 16'hce0;
data_inb = 16'hbf0;
#10;
address_ina = 176;
address_inb = 177;
data_ina = 16'hac2;
data_inb = 16'h0;
#10;
address_ina = 178;
address_inb = 179;
data_ina = 16'h2a7;
data_inb = 16'h751;
#10;
address_ina = 180;
address_inb = 181;
data_ina = 16'h5f1;
data_inb = 16'h747;
#10;
address_ina = 182;
address_inb = 183;
data_ina = 16'h5ba;
data_inb = 16'h9c1;
#10;
address_ina = 184;
address_inb = 185;
data_ina = 16'hc62;
data_inb = 16'h4fa;
#10;
address_ina = 186;
address_inb = 187;
data_ina = 16'h1c4;
data_inb = 16'h653;
#10;
address_ina = 188;
address_inb = 189;
data_ina = 16'h6ae;
data_inb = 16'hac2;
#10;
address_ina = 190;
address_inb = 191;
data_ina = 16'h222;
data_inb = 16'h9c;
#10;
address_ina = 192;
address_inb = 193;
data_ina = 16'h222;
data_inb = 16'h666;
#10;
address_ina = 194;
address_inb = 195;
data_ina = 16'h596;
data_inb = 16'h4ea;
#10;
address_ina = 196;
address_inb = 197;
data_ina = 16'h81a;
data_inb = 16'h482;
#10;
address_ina = 198;
address_inb = 199;
data_ina = 16'h7e6;
data_inb = 16'hbcc;
#10;
address_ina = 200;
address_inb = 201;
data_ina = 16'h95c;
data_inb = 16'h6b5;
#10;
address_ina = 202;
address_inb = 203;
data_ina = 16'h135;
data_inb = 16'h5db;
#10;
address_ina = 204;
address_inb = 205;
data_ina = 16'h9ee;
data_inb = 16'h49f;
#10;
address_ina = 206;
address_inb = 207;
data_ina = 16'h566;
data_inb = 16'h4dd;
#10;
address_ina = 208;
address_inb = 209;
data_ina = 16'hc03;
data_inb = 16'h294;
#10;
address_ina = 210;
address_inb = 211;
data_ina = 16'h148;
data_inb = 16'h911;
#10;
address_ina = 212;
address_inb = 213;
data_ina = 16'h319;
data_inb = 16'hc0;
#10;
address_ina = 214;
address_inb = 215;
data_ina = 16'h764;
data_inb = 16'h148;
#10;
address_ina = 216;
address_inb = 217;
data_ina = 16'ha1c;
data_inb = 16'ha3c;
#10;
address_ina = 218;
address_inb = 219;
data_ina = 16'h13f;
data_inb = 16'h914;
#10;
address_ina = 220;
address_inb = 221;
data_ina = 16'h371;
data_inb = 16'h3e3;
#10;
address_ina = 222;
address_inb = 223;
data_ina = 16'h7b2;
data_inb = 16'h8cd;
#10;
address_ina = 224;
address_inb = 225;
data_ina = 16'h1ad;
data_inb = 16'h6bb;
#10;
address_ina = 226;
address_inb = 227;
data_ina = 16'h65;
data_inb = 16'h25d;
#10;
address_ina = 228;
address_inb = 229;
data_ina = 16'h914;
data_inb = 16'h91e;
#10;
address_ina = 230;
address_inb = 231;
data_ina = 16'h1eb;
data_inb = 16'h6d5;
#10;
address_ina = 232;
address_inb = 233;
data_ina = 16'h973;
data_inb = 16'haef;
#10;
address_ina = 234;
address_inb = 235;
data_ina = 16'h101;
data_inb = 16'h6b;
#10;
address_ina = 236;
address_inb = 237;
data_ina = 16'h132;
data_inb = 16'hab5;
#10;
address_ina = 238;
address_inb = 239;
data_ina = 16'hed;
data_inb = 16'h1a0;
#10;
address_ina = 240;
address_inb = 241;
data_ina = 16'h2d2;
data_inb = 16'h7;
#10;
address_ina = 242;
address_inb = 243;
data_ina = 16'h914;
data_inb = 16'h5a7;
#10;
address_ina = 244;
address_inb = 245;
data_ina = 16'h542;
data_inb = 16'h703;
#10;
address_ina = 246;
address_inb = 247;
data_ina = 16'h19d;
data_inb = 16'h2f2;
#10;
address_ina = 248;
address_inb = 249;
data_ina = 16'h7f6;
data_inb = 16'h69b;
#10;
address_ina = 250;
address_inb = 251;
data_ina = 16'h67d;
data_inb = 16'h650;
#10;
address_ina = 252;
address_inb = 253;
data_ina = 16'h266;
data_inb = 16'h270;
#10;
address_ina = 254;
address_inb = 255;
data_ina = 16'hea;
data_inb = 16'hbb9;
#10;
        wait(init_done);
        #30
        we = 0;
        // Start processing
         
		  #38000

        start = 0;



//        wait (wr_req);
//		  wait (!wr_req);
//		   rd_req = 1;
		  wait(done);
		  #20000
rd_req = 1;
        #70 
		  start = 1;
		 #80 
wait(rd_empty)
rd_req = 0;

$display("Finished the NTT test Number %d",test_num);
////Begin test number #62//////////////
rst = 1;

//#1000
start = 1;
mode = 1; //NTT 0 // INTT 1

// Reset for a few clock cycles

#1000

rst = 0;
test_num = test_num + 1;
#1000
we = 1;
address_ina = 0;
address_inb = 1;
data_ina = 16'hfdee;
data_inb = 16'h55d;
#10;
address_ina = 2;
address_inb = 3;
data_ina = 16'h23f;
data_inb = 16'hfc83;
#10;
address_ina = 4;
address_inb = 5;
data_ina = 16'h66;
data_inb = 16'hfb2f;
#10;
address_ina = 6;
address_inb = 7;
data_ina = 16'hff6c;
data_inb = 16'hfece;
#10;
address_ina = 8;
address_inb = 9;
data_ina = 16'h57b;
data_inb = 16'h330;
#10;
address_ina = 10;
address_inb = 11;
data_ina = 16'hfcde;
data_inb = 16'h16b;
#10;
address_ina = 12;
address_inb = 13;
data_ina = 16'h36;
data_inb = 16'ha8;
#10;
address_ina = 14;
address_inb = 15;
data_ina = 16'h5b;
data_inb = 16'hfa4a;
#10;
address_ina = 16;
address_inb = 17;
data_ina = 16'hfc7b;
data_inb = 16'h40f;
#10;
address_ina = 18;
address_inb = 19;
data_ina = 16'h466;
data_inb = 16'h24d;
#10;
address_ina = 20;
address_inb = 21;
data_ina = 16'h622;
data_inb = 16'hfe4e;
#10;
address_ina = 22;
address_inb = 23;
data_ina = 16'hfe8f;
data_inb = 16'hfacb;
#10;
address_ina = 24;
address_inb = 25;
data_ina = 16'h5cb;
data_inb = 16'hfadc;
#10;
address_ina = 26;
address_inb = 27;
data_ina = 16'h266;
data_inb = 16'h23f;
#10;
address_ina = 28;
address_inb = 29;
data_ina = 16'hfe35;
data_inb = 16'hfe2d;
#10;
address_ina = 30;
address_inb = 31;
data_ina = 16'h66c;
data_inb = 16'hfc48;
#10;
address_ina = 32;
address_inb = 33;
data_ina = 16'h390;
data_inb = 16'hfc56;
#10;
address_ina = 34;
address_inb = 35;
data_ina = 16'hfe35;
data_inb = 16'hfa58;
#10;
address_ina = 36;
address_inb = 37;
data_ina = 16'hfc7f;
data_inb = 16'h32d;
#10;
address_ina = 38;
address_inb = 39;
data_ina = 16'hfc99;
data_inb = 16'hfb4c;
#10;
address_ina = 40;
address_inb = 41;
data_ina = 16'hf98a;
data_inb = 16'h220;
#10;
address_ina = 42;
address_inb = 43;
data_ina = 16'h445;
data_inb = 16'h400;
#10;
address_ina = 44;
address_inb = 45;
data_ina = 16'hfb3b;
data_inb = 16'hfa04;
#10;
address_ina = 46;
address_inb = 47;
data_ina = 16'h363;
data_inb = 16'hfe5e;
#10;
address_ina = 48;
address_inb = 49;
data_ina = 16'h526;
data_inb = 16'hfa30;
#10;
address_ina = 50;
address_inb = 51;
data_ina = 16'h3a7;
data_inb = 16'hfd97;
#10;
address_ina = 52;
address_inb = 53;
data_ina = 16'hfce7;
data_inb = 16'h32;
#10;
address_ina = 54;
address_inb = 55;
data_ina = 16'h1ad;
data_inb = 16'hfa91;
#10;
address_ina = 56;
address_inb = 57;
data_ina = 16'hfbe7;
data_inb = 16'hff04;
#10;
address_ina = 58;
address_inb = 59;
data_ina = 16'h578;
data_inb = 16'hfcee;
#10;
address_ina = 60;
address_inb = 61;
data_ina = 16'hfa3e;
data_inb = 16'h210;
#10;
address_ina = 62;
address_inb = 63;
data_ina = 16'h5a2;
data_inb = 16'h533;
#10;
address_ina = 64;
address_inb = 65;
data_ina = 16'h63c;
data_inb = 16'hfecc;
#10;
address_ina = 66;
address_inb = 67;
data_ina = 16'h2f4;
data_inb = 16'h34e;
#10;
address_ina = 68;
address_inb = 69;
data_ina = 16'h133;
data_inb = 16'hffc8;
#10;
address_ina = 70;
address_inb = 71;
data_ina = 16'hff4f;
data_inb = 16'hf9d7;
#10;
address_ina = 72;
address_inb = 73;
data_ina = 16'hfc63;
data_inb = 16'hfbab;
#10;
address_ina = 74;
address_inb = 75;
data_ina = 16'hfd06;
data_inb = 16'hf9ac;
#10;
address_ina = 76;
address_inb = 77;
data_ina = 16'h2df;
data_inb = 16'h288;
#10;
address_ina = 78;
address_inb = 79;
data_ina = 16'hfb34;
data_inb = 16'h22b;
#10;
address_ina = 80;
address_inb = 81;
data_ina = 16'hfe0d;
data_inb = 16'h18b;
#10;
address_ina = 82;
address_inb = 83;
data_ina = 16'h2be;
data_inb = 16'hee;
#10;
address_ina = 84;
address_inb = 85;
data_ina = 16'hfa74;
data_inb = 16'hfe0d;
#10;
address_ina = 86;
address_inb = 87;
data_ina = 16'h1c7;
data_inb = 16'h171;
#10;
address_ina = 88;
address_inb = 89;
data_ina = 16'haf;
data_inb = 16'hb2;
#10;
address_ina = 90;
address_inb = 91;
data_ina = 16'hfe11;
data_inb = 16'h17d;
#10;
address_ina = 92;
address_inb = 93;
data_ina = 16'hfa81;
data_inb = 16'hfece;
#10;
address_ina = 94;
address_inb = 95;
data_ina = 16'h4f3;
data_inb = 16'h61c;
#10;
address_ina = 96;
address_inb = 97;
data_ina = 16'hfa46;
data_inb = 16'h321;
#10;
address_ina = 98;
address_inb = 99;
data_ina = 16'h3f3;
data_inb = 16'h508;
#10;
address_ina = 100;
address_inb = 101;
data_ina = 16'ha0;
data_inb = 16'h53d;
#10;
address_ina = 102;
address_inb = 103;
data_ina = 16'h410;
data_inb = 16'hfc9c;
#10;
address_ina = 104;
address_inb = 105;
data_ina = 16'h484;
data_inb = 16'hf9ff;
#10;
address_ina = 106;
address_inb = 107;
data_ina = 16'hffe1;
data_inb = 16'hfb59;
#10;
address_ina = 108;
address_inb = 109;
data_ina = 16'hfb7a;
data_inb = 16'hfd94;
#10;
address_ina = 110;
address_inb = 111;
data_ina = 16'h482;
data_inb = 16'hfdd6;
#10;
address_ina = 112;
address_inb = 113;
data_ina = 16'h38f;
data_inb = 16'h2d5;
#10;
address_ina = 114;
address_inb = 115;
data_ina = 16'h61e;
data_inb = 16'hfe89;
#10;
address_ina = 116;
address_inb = 117;
data_ina = 16'hffeb;
data_inb = 16'hfc67;
#10;
address_ina = 118;
address_inb = 119;
data_ina = 16'h615;
data_inb = 16'hfb94;
#10;
address_ina = 120;
address_inb = 121;
data_ina = 16'hfdbc;
data_inb = 16'hfbbb;
#10;
address_ina = 122;
address_inb = 123;
data_ina = 16'hfa81;
data_inb = 16'h52d;
#10;
address_ina = 124;
address_inb = 125;
data_ina = 16'hfe36;
data_inb = 16'h2c7;
#10;
address_ina = 126;
address_inb = 127;
data_ina = 16'h5f7;
data_inb = 16'h3a1;
#10;
address_ina = 128;
address_inb = 129;
data_ina = 16'h4c4;
data_inb = 16'h176;
#10;
address_ina = 130;
address_inb = 131;
data_ina = 16'h31a;
data_inb = 16'h86;
#10;
address_ina = 132;
address_inb = 133;
data_ina = 16'hfffc;
data_inb = 16'h415;
#10;
address_ina = 134;
address_inb = 135;
data_ina = 16'hfe79;
data_inb = 16'h21c;
#10;
address_ina = 136;
address_inb = 137;
data_ina = 16'h20a;
data_inb = 16'hb8;
#10;
address_ina = 138;
address_inb = 139;
data_ina = 16'hfef3;
data_inb = 16'hfa8e;
#10;
address_ina = 140;
address_inb = 141;
data_ina = 16'hfba5;
data_inb = 16'h11c;
#10;
address_ina = 142;
address_inb = 143;
data_ina = 16'hfdd7;
data_inb = 16'h556;
#10;
address_ina = 144;
address_inb = 145;
data_ina = 16'hfeef;
data_inb = 16'hfb6c;
#10;
address_ina = 146;
address_inb = 147;
data_ina = 16'h4e5;
data_inb = 16'hfeb9;
#10;
address_ina = 148;
address_inb = 149;
data_ina = 16'h489;
data_inb = 16'h58;
#10;
address_ina = 150;
address_inb = 151;
data_ina = 16'h638;
data_inb = 16'ha6;
#10;
address_ina = 152;
address_inb = 153;
data_ina = 16'hfeaa;
data_inb = 16'h566;
#10;
address_ina = 154;
address_inb = 155;
data_ina = 16'h237;
data_inb = 16'hfb38;
#10;
address_ina = 156;
address_inb = 157;
data_ina = 16'haf;
data_inb = 16'h94;
#10;
address_ina = 158;
address_inb = 159;
data_ina = 16'h5b3;
data_inb = 16'he1;
#10;
address_ina = 160;
address_inb = 161;
data_ina = 16'h1f5;
data_inb = 16'h252;
#10;
address_ina = 162;
address_inb = 163;
data_ina = 16'hf9ec;
data_inb = 16'h35f;
#10;
address_ina = 164;
address_inb = 165;
data_ina = 16'hfe1e;
data_inb = 16'h69;
#10;
address_ina = 166;
address_inb = 167;
data_ina = 16'h2d3;
data_inb = 16'h364;
#10;
address_ina = 168;
address_inb = 169;
data_ina = 16'hfae9;
data_inb = 16'h19;
#10;
address_ina = 170;
address_inb = 171;
data_ina = 16'hfb6a;
data_inb = 16'h20a;
#10;
address_ina = 172;
address_inb = 173;
data_ina = 16'hfff1;
data_inb = 16'h126;
#10;
address_ina = 174;
address_inb = 175;
data_ina = 16'h309;
data_inb = 16'hfa52;
#10;
address_ina = 176;
address_inb = 177;
data_ina = 16'h444;
data_inb = 16'hfd12;
#10;
address_ina = 178;
address_inb = 179;
data_ina = 16'h195;
data_inb = 16'hc1;
#10;
address_ina = 180;
address_inb = 181;
data_ina = 16'h3ad;
data_inb = 16'h4e8;
#10;
address_ina = 182;
address_inb = 183;
data_ina = 16'hf9dd;
data_inb = 16'hff7d;
#10;
address_ina = 184;
address_inb = 185;
data_ina = 16'hfbac;
data_inb = 16'hff98;
#10;
address_ina = 186;
address_inb = 187;
data_ina = 16'h2f4;
data_inb = 16'h2d1;
#10;
address_ina = 188;
address_inb = 189;
data_ina = 16'hf9ac;
data_inb = 16'hfb09;
#10;
address_ina = 190;
address_inb = 191;
data_ina = 16'hfa22;
data_inb = 16'hff48;
#10;
address_ina = 192;
address_inb = 193;
data_ina = 16'hfdba;
data_inb = 16'h292;
#10;
address_ina = 194;
address_inb = 195;
data_ina = 16'hfc29;
data_inb = 16'hfcba;
#10;
address_ina = 196;
address_inb = 197;
data_ina = 16'h2ee;
data_inb = 16'h443;
#10;
address_ina = 198;
address_inb = 199;
data_ina = 16'hfb31;
data_inb = 16'hfacc;
#10;
address_ina = 200;
address_inb = 201;
data_ina = 16'h31d;
data_inb = 16'hfb28;
#10;
address_ina = 202;
address_inb = 203;
data_ina = 16'hfbfa;
data_inb = 16'hfe7d;
#10;
address_ina = 204;
address_inb = 205;
data_ina = 16'hfdee;
data_inb = 16'hfa43;
#10;
address_ina = 206;
address_inb = 207;
data_ina = 16'hfb8f;
data_inb = 16'hf9ae;
#10;
address_ina = 208;
address_inb = 209;
data_ina = 16'h5de;
data_inb = 16'hff15;
#10;
address_ina = 210;
address_inb = 211;
data_ina = 16'h433;
data_inb = 16'hfbe0;
#10;
address_ina = 212;
address_inb = 213;
data_ina = 16'h339;
data_inb = 16'h548;
#10;
address_ina = 214;
address_inb = 215;
data_ina = 16'h3ec;
data_inb = 16'h138;
#10;
address_ina = 216;
address_inb = 217;
data_ina = 16'h453;
data_inb = 16'hf984;
#10;
address_ina = 218;
address_inb = 219;
data_ina = 16'h3a4;
data_inb = 16'h267;
#10;
address_ina = 220;
address_inb = 221;
data_ina = 16'hfdc6;
data_inb = 16'hfc7d;
#10;
address_ina = 222;
address_inb = 223;
data_ina = 16'hfb8e;
data_inb = 16'h112;
#10;
address_ina = 224;
address_inb = 225;
data_ina = 16'he1;
data_inb = 16'hfb6e;
#10;
address_ina = 226;
address_inb = 227;
data_ina = 16'h408;
data_inb = 16'hfd5f;
#10;
address_ina = 228;
address_inb = 229;
data_ina = 16'h212;
data_inb = 16'h157;
#10;
address_ina = 230;
address_inb = 231;
data_ina = 16'hfe96;
data_inb = 16'h97;
#10;
address_ina = 232;
address_inb = 233;
data_ina = 16'h25b;
data_inb = 16'hfc19;
#10;
address_ina = 234;
address_inb = 235;
data_ina = 16'hfe43;
data_inb = 16'h340;
#10;
address_ina = 236;
address_inb = 237;
data_ina = 16'hf9a5;
data_inb = 16'h1fe;
#10;
address_ina = 238;
address_inb = 239;
data_ina = 16'h29d;
data_inb = 16'hfc8b;
#10;
address_ina = 240;
address_inb = 241;
data_ina = 16'h24e;
data_inb = 16'h2f6;
#10;
address_ina = 242;
address_inb = 243;
data_ina = 16'hffef;
data_inb = 16'hff8b;
#10;
address_ina = 244;
address_inb = 245;
data_ina = 16'h3e8;
data_inb = 16'h15d;
#10;
address_ina = 246;
address_inb = 247;
data_ina = 16'hfb38;
data_inb = 16'hff68;
#10;
address_ina = 248;
address_inb = 249;
data_ina = 16'hfd44;
data_inb = 16'hfd9f;
#10;
address_ina = 250;
address_inb = 251;
data_ina = 16'hfda7;
data_inb = 16'h283;
#10;
address_ina = 252;
address_inb = 253;
data_ina = 16'hfe96;
data_inb = 16'h2a;
#10;
address_ina = 254;
address_inb = 255;
data_ina = 16'h19d;
data_inb = 16'hfffb;
#10;
        wait(init_done);
        #30
        we = 0;
        // Start processing
         
		  #38000

        start = 0;



//        wait (wr_req);
//		  wait (!wr_req);
//		   rd_req = 1;
		  wait(done);
		  #20000
rd_req = 1;
        #70 
		  start = 1;
		 #80 
wait(rd_empty)
rd_req = 0;

$display("Finished the NTT test Number %d",test_num);
////Begin test number #63//////////////
rst = 1;

//#1000
start = 1;
mode = 0; //NTT 0 // INTT 1

// Reset for a few clock cycles

#1000

rst = 0;
test_num = test_num + 1;
#1000
we = 1;
address_ina = 0;
address_inb = 1;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 2;
address_inb = 3;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 4;
address_inb = 5;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 6;
address_inb = 7;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 8;
address_inb = 9;
data_ina = 16'h2;
data_inb = 16'h0;
#10;
address_ina = 10;
address_inb = 11;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 12;
address_inb = 13;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 14;
address_inb = 15;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 16;
address_inb = 17;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 18;
address_inb = 19;
data_ina = 16'hfffd;
data_inb = 16'h1;
#10;
address_ina = 20;
address_inb = 21;
data_ina = 16'h1;
data_inb = 16'h2;
#10;
address_ina = 22;
address_inb = 23;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 24;
address_inb = 25;
data_ina = 16'h1;
data_inb = 16'h2;
#10;
address_ina = 26;
address_inb = 27;
data_ina = 16'h2;
data_inb = 16'h1;
#10;
address_ina = 28;
address_inb = 29;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 30;
address_inb = 31;
data_ina = 16'h2;
data_inb = 16'h2;
#10;
address_ina = 32;
address_inb = 33;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 34;
address_inb = 35;
data_ina = 16'h0;
data_inb = 16'hfffe;
#10;
address_ina = 36;
address_inb = 37;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 38;
address_inb = 39;
data_ina = 16'hfffe;
data_inb = 16'hffff;
#10;
address_ina = 40;
address_inb = 41;
data_ina = 16'h0;
data_inb = 16'hfffd;
#10;
address_ina = 42;
address_inb = 43;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 44;
address_inb = 45;
data_ina = 16'hfffe;
data_inb = 16'hffff;
#10;
address_ina = 46;
address_inb = 47;
data_ina = 16'h3;
data_inb = 16'hfffd;
#10;
address_ina = 48;
address_inb = 49;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 50;
address_inb = 51;
data_ina = 16'h3;
data_inb = 16'h0;
#10;
address_ina = 52;
address_inb = 53;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 54;
address_inb = 55;
data_ina = 16'hfffd;
data_inb = 16'h1;
#10;
address_ina = 56;
address_inb = 57;
data_ina = 16'hffff;
data_inb = 16'hfffe;
#10;
address_ina = 58;
address_inb = 59;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 60;
address_inb = 61;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 62;
address_inb = 63;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 64;
address_inb = 65;
data_ina = 16'hfffe;
data_inb = 16'h1;
#10;
address_ina = 66;
address_inb = 67;
data_ina = 16'h2;
data_inb = 16'h2;
#10;
address_ina = 68;
address_inb = 69;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 70;
address_inb = 71;
data_ina = 16'hfffe;
data_inb = 16'hfffd;
#10;
address_ina = 72;
address_inb = 73;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 74;
address_inb = 75;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 76;
address_inb = 77;
data_ina = 16'hffff;
data_inb = 16'h2;
#10;
address_ina = 78;
address_inb = 79;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 80;
address_inb = 81;
data_ina = 16'h0;
data_inb = 16'hfffe;
#10;
address_ina = 82;
address_inb = 83;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 84;
address_inb = 85;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 86;
address_inb = 87;
data_ina = 16'h2;
data_inb = 16'h0;
#10;
address_ina = 88;
address_inb = 89;
data_ina = 16'h3;
data_inb = 16'hffff;
#10;
address_ina = 90;
address_inb = 91;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 92;
address_inb = 93;
data_ina = 16'hffff;
data_inb = 16'hfffd;
#10;
address_ina = 94;
address_inb = 95;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 96;
address_inb = 97;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 98;
address_inb = 99;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 100;
address_inb = 101;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 102;
address_inb = 103;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 104;
address_inb = 105;
data_ina = 16'h2;
data_inb = 16'h1;
#10;
address_ina = 106;
address_inb = 107;
data_ina = 16'hffff;
data_inb = 16'h2;
#10;
address_ina = 108;
address_inb = 109;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 110;
address_inb = 111;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 112;
address_inb = 113;
data_ina = 16'h0;
data_inb = 16'h3;
#10;
address_ina = 114;
address_inb = 115;
data_ina = 16'hfffe;
data_inb = 16'h1;
#10;
address_ina = 116;
address_inb = 117;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 118;
address_inb = 119;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 120;
address_inb = 121;
data_ina = 16'hfffe;
data_inb = 16'hfffe;
#10;
address_ina = 122;
address_inb = 123;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 124;
address_inb = 125;
data_ina = 16'h0;
data_inb = 16'hfffe;
#10;
address_ina = 126;
address_inb = 127;
data_ina = 16'h2;
data_inb = 16'hfffe;
#10;
address_ina = 128;
address_inb = 129;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 130;
address_inb = 131;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 132;
address_inb = 133;
data_ina = 16'hffff;
data_inb = 16'hfffe;
#10;
address_ina = 134;
address_inb = 135;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 136;
address_inb = 137;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 138;
address_inb = 139;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 140;
address_inb = 141;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 142;
address_inb = 143;
data_ina = 16'h2;
data_inb = 16'h1;
#10;
address_ina = 144;
address_inb = 145;
data_ina = 16'hffff;
data_inb = 16'hfffe;
#10;
address_ina = 146;
address_inb = 147;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 148;
address_inb = 149;
data_ina = 16'h0;
data_inb = 16'hfffe;
#10;
address_ina = 150;
address_inb = 151;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 152;
address_inb = 153;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 154;
address_inb = 155;
data_ina = 16'hfffd;
data_inb = 16'h1;
#10;
address_ina = 156;
address_inb = 157;
data_ina = 16'h2;
data_inb = 16'hffff;
#10;
address_ina = 158;
address_inb = 159;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 160;
address_inb = 161;
data_ina = 16'h3;
data_inb = 16'h0;
#10;
address_ina = 162;
address_inb = 163;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 164;
address_inb = 165;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 166;
address_inb = 167;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 168;
address_inb = 169;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 170;
address_inb = 171;
data_ina = 16'h1;
data_inb = 16'h3;
#10;
address_ina = 172;
address_inb = 173;
data_ina = 16'h0;
data_inb = 16'h2;
#10;
address_ina = 174;
address_inb = 175;
data_ina = 16'h1;
data_inb = 16'h3;
#10;
address_ina = 176;
address_inb = 177;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 178;
address_inb = 179;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 180;
address_inb = 181;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 182;
address_inb = 183;
data_ina = 16'hfffd;
data_inb = 16'h0;
#10;
address_ina = 184;
address_inb = 185;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 186;
address_inb = 187;
data_ina = 16'h3;
data_inb = 16'hffff;
#10;
address_ina = 188;
address_inb = 189;
data_ina = 16'hffff;
data_inb = 16'hfffe;
#10;
address_ina = 190;
address_inb = 191;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 192;
address_inb = 193;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 194;
address_inb = 195;
data_ina = 16'h2;
data_inb = 16'h0;
#10;
address_ina = 196;
address_inb = 197;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 198;
address_inb = 199;
data_ina = 16'h0;
data_inb = 16'h2;
#10;
address_ina = 200;
address_inb = 201;
data_ina = 16'hfffe;
data_inb = 16'h0;
#10;
address_ina = 202;
address_inb = 203;
data_ina = 16'h2;
data_inb = 16'h0;
#10;
address_ina = 204;
address_inb = 205;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 206;
address_inb = 207;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 208;
address_inb = 209;
data_ina = 16'h1;
data_inb = 16'h2;
#10;
address_ina = 210;
address_inb = 211;
data_ina = 16'hffff;
data_inb = 16'h2;
#10;
address_ina = 212;
address_inb = 213;
data_ina = 16'hfffe;
data_inb = 16'h1;
#10;
address_ina = 214;
address_inb = 215;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 216;
address_inb = 217;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 218;
address_inb = 219;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 220;
address_inb = 221;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 222;
address_inb = 223;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 224;
address_inb = 225;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 226;
address_inb = 227;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 228;
address_inb = 229;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 230;
address_inb = 231;
data_ina = 16'h1;
data_inb = 16'hfffd;
#10;
address_ina = 232;
address_inb = 233;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 234;
address_inb = 235;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 236;
address_inb = 237;
data_ina = 16'hfffe;
data_inb = 16'h1;
#10;
address_ina = 238;
address_inb = 239;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 240;
address_inb = 241;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 242;
address_inb = 243;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 244;
address_inb = 245;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 246;
address_inb = 247;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 248;
address_inb = 249;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 250;
address_inb = 251;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 252;
address_inb = 253;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 254;
address_inb = 255;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
        wait(init_done);
        #30
        we = 0;
        // Start processing
         
		  #38000

        start = 0;



//        wait (wr_req);
//		  wait (!wr_req);
//		   rd_req = 1;
		  wait(done);
		  #20000
rd_req = 1;
        #70 
		  start = 1;
		 #80 
wait(rd_empty)
rd_req = 0;

$display("Finished the NTT test Number %d",test_num);
////Begin test number #64//////////////
rst = 1;

//#1000
start = 1;
mode = 0; //NTT 0 // INTT 1

// Reset for a few clock cycles

#1000

rst = 0;
test_num = test_num + 1;
#1000
we = 1;
address_ina = 0;
address_inb = 1;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 2;
address_inb = 3;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 4;
address_inb = 5;
data_ina = 16'hfffe;
data_inb = 16'h1;
#10;
address_ina = 6;
address_inb = 7;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 8;
address_inb = 9;
data_ina = 16'h3;
data_inb = 16'h0;
#10;
address_ina = 10;
address_inb = 11;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 12;
address_inb = 13;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 14;
address_inb = 15;
data_ina = 16'hffff;
data_inb = 16'hfffe;
#10;
address_ina = 16;
address_inb = 17;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 18;
address_inb = 19;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 20;
address_inb = 21;
data_ina = 16'hfffe;
data_inb = 16'h0;
#10;
address_ina = 22;
address_inb = 23;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 24;
address_inb = 25;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 26;
address_inb = 27;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 28;
address_inb = 29;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 30;
address_inb = 31;
data_ina = 16'h1;
data_inb = 16'h3;
#10;
address_ina = 32;
address_inb = 33;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 34;
address_inb = 35;
data_ina = 16'hfffe;
data_inb = 16'h1;
#10;
address_ina = 36;
address_inb = 37;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 38;
address_inb = 39;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 40;
address_inb = 41;
data_ina = 16'h0;
data_inb = 16'hfffe;
#10;
address_ina = 42;
address_inb = 43;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 44;
address_inb = 45;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 46;
address_inb = 47;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 48;
address_inb = 49;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 50;
address_inb = 51;
data_ina = 16'hfffe;
data_inb = 16'hffff;
#10;
address_ina = 52;
address_inb = 53;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 54;
address_inb = 55;
data_ina = 16'h1;
data_inb = 16'hfffd;
#10;
address_ina = 56;
address_inb = 57;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 58;
address_inb = 59;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 60;
address_inb = 61;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 62;
address_inb = 63;
data_ina = 16'hfffe;
data_inb = 16'h0;
#10;
address_ina = 64;
address_inb = 65;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 66;
address_inb = 67;
data_ina = 16'hffff;
data_inb = 16'hfffe;
#10;
address_ina = 68;
address_inb = 69;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 70;
address_inb = 71;
data_ina = 16'h0;
data_inb = 16'h2;
#10;
address_ina = 72;
address_inb = 73;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 74;
address_inb = 75;
data_ina = 16'h1;
data_inb = 16'hfffe;
#10;
address_ina = 76;
address_inb = 77;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 78;
address_inb = 79;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 80;
address_inb = 81;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 82;
address_inb = 83;
data_ina = 16'hffff;
data_inb = 16'h2;
#10;
address_ina = 84;
address_inb = 85;
data_ina = 16'h2;
data_inb = 16'hfffd;
#10;
address_ina = 86;
address_inb = 87;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 88;
address_inb = 89;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 90;
address_inb = 91;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 92;
address_inb = 93;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 94;
address_inb = 95;
data_ina = 16'h1;
data_inb = 16'hfffe;
#10;
address_ina = 96;
address_inb = 97;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 98;
address_inb = 99;
data_ina = 16'h0;
data_inb = 16'h2;
#10;
address_ina = 100;
address_inb = 101;
data_ina = 16'hfffe;
data_inb = 16'hffff;
#10;
address_ina = 102;
address_inb = 103;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 104;
address_inb = 105;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 106;
address_inb = 107;
data_ina = 16'h2;
data_inb = 16'hffff;
#10;
address_ina = 108;
address_inb = 109;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 110;
address_inb = 111;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 112;
address_inb = 113;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 114;
address_inb = 115;
data_ina = 16'h2;
data_inb = 16'h1;
#10;
address_ina = 116;
address_inb = 117;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 118;
address_inb = 119;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 120;
address_inb = 121;
data_ina = 16'hfffe;
data_inb = 16'h1;
#10;
address_ina = 122;
address_inb = 123;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 124;
address_inb = 125;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 126;
address_inb = 127;
data_ina = 16'h2;
data_inb = 16'h0;
#10;
address_ina = 128;
address_inb = 129;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 130;
address_inb = 131;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 132;
address_inb = 133;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 134;
address_inb = 135;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 136;
address_inb = 137;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 138;
address_inb = 139;
data_ina = 16'hffff;
data_inb = 16'h2;
#10;
address_ina = 140;
address_inb = 141;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 142;
address_inb = 143;
data_ina = 16'h1;
data_inb = 16'hfffe;
#10;
address_ina = 144;
address_inb = 145;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 146;
address_inb = 147;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 148;
address_inb = 149;
data_ina = 16'h2;
data_inb = 16'h2;
#10;
address_ina = 150;
address_inb = 151;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 152;
address_inb = 153;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 154;
address_inb = 155;
data_ina = 16'hffff;
data_inb = 16'h2;
#10;
address_ina = 156;
address_inb = 157;
data_ina = 16'hfffe;
data_inb = 16'hffff;
#10;
address_ina = 158;
address_inb = 159;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 160;
address_inb = 161;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 162;
address_inb = 163;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 164;
address_inb = 165;
data_ina = 16'hfffd;
data_inb = 16'hffff;
#10;
address_ina = 166;
address_inb = 167;
data_ina = 16'hfffe;
data_inb = 16'h0;
#10;
address_ina = 168;
address_inb = 169;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 170;
address_inb = 171;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 172;
address_inb = 173;
data_ina = 16'h1;
data_inb = 16'hfffe;
#10;
address_ina = 174;
address_inb = 175;
data_ina = 16'hfffe;
data_inb = 16'h1;
#10;
address_ina = 176;
address_inb = 177;
data_ina = 16'hffff;
data_inb = 16'h2;
#10;
address_ina = 178;
address_inb = 179;
data_ina = 16'hfffe;
data_inb = 16'h0;
#10;
address_ina = 180;
address_inb = 181;
data_ina = 16'h1;
data_inb = 16'h2;
#10;
address_ina = 182;
address_inb = 183;
data_ina = 16'hffff;
data_inb = 16'h3;
#10;
address_ina = 184;
address_inb = 185;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 186;
address_inb = 187;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 188;
address_inb = 189;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 190;
address_inb = 191;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 192;
address_inb = 193;
data_ina = 16'hffff;
data_inb = 16'hfffe;
#10;
address_ina = 194;
address_inb = 195;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 196;
address_inb = 197;
data_ina = 16'h0;
data_inb = 16'hfffe;
#10;
address_ina = 198;
address_inb = 199;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 200;
address_inb = 201;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 202;
address_inb = 203;
data_ina = 16'h2;
data_inb = 16'h0;
#10;
address_ina = 204;
address_inb = 205;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 206;
address_inb = 207;
data_ina = 16'hfffd;
data_inb = 16'hfffe;
#10;
address_ina = 208;
address_inb = 209;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 210;
address_inb = 211;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 212;
address_inb = 213;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 214;
address_inb = 215;
data_ina = 16'h0;
data_inb = 16'h2;
#10;
address_ina = 216;
address_inb = 217;
data_ina = 16'h2;
data_inb = 16'h1;
#10;
address_ina = 218;
address_inb = 219;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 220;
address_inb = 221;
data_ina = 16'h3;
data_inb = 16'h1;
#10;
address_ina = 222;
address_inb = 223;
data_ina = 16'h2;
data_inb = 16'hffff;
#10;
address_ina = 224;
address_inb = 225;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 226;
address_inb = 227;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 228;
address_inb = 229;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 230;
address_inb = 231;
data_ina = 16'h2;
data_inb = 16'h1;
#10;
address_ina = 232;
address_inb = 233;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 234;
address_inb = 235;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 236;
address_inb = 237;
data_ina = 16'h0;
data_inb = 16'hfffe;
#10;
address_ina = 238;
address_inb = 239;
data_ina = 16'h0;
data_inb = 16'hfffe;
#10;
address_ina = 240;
address_inb = 241;
data_ina = 16'hfffe;
data_inb = 16'hfffe;
#10;
address_ina = 242;
address_inb = 243;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 244;
address_inb = 245;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 246;
address_inb = 247;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 248;
address_inb = 249;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 250;
address_inb = 251;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 252;
address_inb = 253;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 254;
address_inb = 255;
data_ina = 16'h1;
data_inb = 16'h2;
#10;
        wait(init_done);
        #30
        we = 0;
        // Start processing
         
		  #38000

        start = 0;



//        wait (wr_req);
//		  wait (!wr_req);
//		   rd_req = 1;
		  wait(done);
		  #20000
rd_req = 1;
        #70 
		  start = 1;
		 #80 
wait(rd_empty)
rd_req = 0;

$display("Finished the NTT test Number %d",test_num);
////Begin test number #65//////////////
rst = 1;

//#1000
start = 1;
mode = 1; //NTT 0 // INTT 1

// Reset for a few clock cycles

#1000

rst = 0;
test_num = test_num + 1;
#1000
we = 1;
address_ina = 0;
address_inb = 1;
data_ina = 16'hfc36;
data_inb = 16'ha5;
#10;
address_ina = 2;
address_inb = 3;
data_ina = 16'h4b3;
data_inb = 16'h22b;
#10;
address_ina = 4;
address_inb = 5;
data_ina = 16'hfb68;
data_inb = 16'hc4;
#10;
address_ina = 6;
address_inb = 7;
data_ina = 16'hfb62;
data_inb = 16'hfb88;
#10;
address_ina = 8;
address_inb = 9;
data_ina = 16'hf0;
data_inb = 16'hfa50;
#10;
address_ina = 10;
address_inb = 11;
data_ina = 16'hfb45;
data_inb = 16'h17;
#10;
address_ina = 12;
address_inb = 13;
data_ina = 16'h11c;
data_inb = 16'hc0;
#10;
address_ina = 14;
address_inb = 15;
data_ina = 16'hfa7e;
data_inb = 16'hfdd0;
#10;
address_ina = 16;
address_inb = 17;
data_ina = 16'hff51;
data_inb = 16'h468;
#10;
address_ina = 18;
address_inb = 19;
data_ina = 16'hfd2a;
data_inb = 16'h30b;
#10;
address_ina = 20;
address_inb = 21;
data_ina = 16'h412;
data_inb = 16'hfeb3;
#10;
address_ina = 22;
address_inb = 23;
data_ina = 16'h50b;
data_inb = 16'hfbe6;
#10;
address_ina = 24;
address_inb = 25;
data_ina = 16'hfb43;
data_inb = 16'h3ee;
#10;
address_ina = 26;
address_inb = 27;
data_ina = 16'h196;
data_inb = 16'hff28;
#10;
address_ina = 28;
address_inb = 29;
data_ina = 16'hfe59;
data_inb = 16'hfa6d;
#10;
address_ina = 30;
address_inb = 31;
data_ina = 16'h3b5;
data_inb = 16'h593;
#10;
address_ina = 32;
address_inb = 33;
data_ina = 16'hfb2e;
data_inb = 16'hfeb4;
#10;
address_ina = 34;
address_inb = 35;
data_ina = 16'h475;
data_inb = 16'h386;
#10;
address_ina = 36;
address_inb = 37;
data_ina = 16'hfab1;
data_inb = 16'h3f4;
#10;
address_ina = 38;
address_inb = 39;
data_ina = 16'hfe17;
data_inb = 16'hfc5e;
#10;
address_ina = 40;
address_inb = 41;
data_ina = 16'hfe8c;
data_inb = 16'hfcd6;
#10;
address_ina = 42;
address_inb = 43;
data_ina = 16'hfa34;
data_inb = 16'hfbc8;
#10;
address_ina = 44;
address_inb = 45;
data_ina = 16'h3d9;
data_inb = 16'h40b;
#10;
address_ina = 46;
address_inb = 47;
data_ina = 16'hf9ed;
data_inb = 16'h32;
#10;
address_ina = 48;
address_inb = 49;
data_ina = 16'h282;
data_inb = 16'h52;
#10;
address_ina = 50;
address_inb = 51;
data_ina = 16'hf9c5;
data_inb = 16'h4bb;
#10;
address_ina = 52;
address_inb = 53;
data_ina = 16'hfd1d;
data_inb = 16'h7a;
#10;
address_ina = 54;
address_inb = 55;
data_ina = 16'hfa8e;
data_inb = 16'hff38;
#10;
address_ina = 56;
address_inb = 57;
data_ina = 16'h22;
data_inb = 16'hfc59;
#10;
address_ina = 58;
address_inb = 59;
data_ina = 16'h51c;
data_inb = 16'h581;
#10;
address_ina = 60;
address_inb = 61;
data_ina = 16'hfb57;
data_inb = 16'h542;
#10;
address_ina = 62;
address_inb = 63;
data_ina = 16'h608;
data_inb = 16'h573;
#10;
address_ina = 64;
address_inb = 65;
data_ina = 16'h535;
data_inb = 16'hff9e;
#10;
address_ina = 66;
address_inb = 67;
data_ina = 16'hfe9a;
data_inb = 16'hfa3d;
#10;
address_ina = 68;
address_inb = 69;
data_ina = 16'h2a;
data_inb = 16'h671;
#10;
address_ina = 70;
address_inb = 71;
data_ina = 16'hffc4;
data_inb = 16'h59a;
#10;
address_ina = 72;
address_inb = 73;
data_ina = 16'hfb05;
data_inb = 16'hf995;
#10;
address_ina = 74;
address_inb = 75;
data_ina = 16'h352;
data_inb = 16'hfc88;
#10;
address_ina = 76;
address_inb = 77;
data_ina = 16'h642;
data_inb = 16'hfd4c;
#10;
address_ina = 78;
address_inb = 79;
data_ina = 16'hfdea;
data_inb = 16'hffb2;
#10;
address_ina = 80;
address_inb = 81;
data_ina = 16'hfb18;
data_inb = 16'hfd53;
#10;
address_ina = 82;
address_inb = 83;
data_ina = 16'hfaf7;
data_inb = 16'h5f6;
#10;
address_ina = 84;
address_inb = 85;
data_ina = 16'h67a;
data_inb = 16'hff9c;
#10;
address_ina = 86;
address_inb = 87;
data_ina = 16'h566;
data_inb = 16'h302;
#10;
address_ina = 88;
address_inb = 89;
data_ina = 16'h2fa;
data_inb = 16'h4e2;
#10;
address_ina = 90;
address_inb = 91;
data_ina = 16'h411;
data_inb = 16'hfbe2;
#10;
address_ina = 92;
address_inb = 93;
data_ina = 16'hfe68;
data_inb = 16'hf9a7;
#10;
address_ina = 94;
address_inb = 95;
data_ina = 16'hfd7b;
data_inb = 16'h32b;
#10;
address_ina = 96;
address_inb = 97;
data_ina = 16'h7f;
data_inb = 16'hfdbc;
#10;
address_ina = 98;
address_inb = 99;
data_ina = 16'hfc59;
data_inb = 16'hfb21;
#10;
address_ina = 100;
address_inb = 101;
data_ina = 16'hff3c;
data_inb = 16'h2a7;
#10;
address_ina = 102;
address_inb = 103;
data_ina = 16'h3f2;
data_inb = 16'h623;
#10;
address_ina = 104;
address_inb = 105;
data_ina = 16'h56e;
data_inb = 16'hfe29;
#10;
address_ina = 106;
address_inb = 107;
data_ina = 16'h57;
data_inb = 16'hfd15;
#10;
address_ina = 108;
address_inb = 109;
data_ina = 16'hfee6;
data_inb = 16'hff88;
#10;
address_ina = 110;
address_inb = 111;
data_ina = 16'h518;
data_inb = 16'h627;
#10;
address_ina = 112;
address_inb = 113;
data_ina = 16'h435;
data_inb = 16'h302;
#10;
address_ina = 114;
address_inb = 115;
data_ina = 16'hfb00;
data_inb = 16'h298;
#10;
address_ina = 116;
address_inb = 117;
data_ina = 16'hfb3f;
data_inb = 16'hf9eb;
#10;
address_ina = 118;
address_inb = 119;
data_ina = 16'h623;
data_inb = 16'hfb86;
#10;
address_ina = 120;
address_inb = 121;
data_ina = 16'hf9dc;
data_inb = 16'hf997;
#10;
address_ina = 122;
address_inb = 123;
data_ina = 16'hfacf;
data_inb = 16'hffef;
#10;
address_ina = 124;
address_inb = 125;
data_ina = 16'hfe6f;
data_inb = 16'h1e5;
#10;
address_ina = 126;
address_inb = 127;
data_ina = 16'h52a;
data_inb = 16'hfbc0;
#10;
address_ina = 128;
address_inb = 129;
data_ina = 16'h89;
data_inb = 16'h455;
#10;
address_ina = 130;
address_inb = 131;
data_ina = 16'hfa22;
data_inb = 16'hff5b;
#10;
address_ina = 132;
address_inb = 133;
data_ina = 16'h269;
data_inb = 16'hfce6;
#10;
address_ina = 134;
address_inb = 135;
data_ina = 16'hff5e;
data_inb = 16'hfd1c;
#10;
address_ina = 136;
address_inb = 137;
data_ina = 16'hfedd;
data_inb = 16'hffae;
#10;
address_ina = 138;
address_inb = 139;
data_ina = 16'h667;
data_inb = 16'h3a3;
#10;
address_ina = 140;
address_inb = 141;
data_ina = 16'h4dd;
data_inb = 16'h16f;
#10;
address_ina = 142;
address_inb = 143;
data_ina = 16'h535;
data_inb = 16'h344;
#10;
address_ina = 144;
address_inb = 145;
data_ina = 16'hff25;
data_inb = 16'h159;
#10;
address_ina = 146;
address_inb = 147;
data_ina = 16'hf9b7;
data_inb = 16'hfe91;
#10;
address_ina = 148;
address_inb = 149;
data_ina = 16'h4aa;
data_inb = 16'hfa15;
#10;
address_ina = 150;
address_inb = 151;
data_ina = 16'hfa82;
data_inb = 16'h536;
#10;
address_ina = 152;
address_inb = 153;
data_ina = 16'hffe7;
data_inb = 16'h3b2;
#10;
address_ina = 154;
address_inb = 155;
data_ina = 16'h85;
data_inb = 16'h183;
#10;
address_ina = 156;
address_inb = 157;
data_ina = 16'hfa43;
data_inb = 16'h242;
#10;
address_ina = 158;
address_inb = 159;
data_ina = 16'hfc4a;
data_inb = 16'hfb26;
#10;
address_ina = 160;
address_inb = 161;
data_ina = 16'hfec8;
data_inb = 16'hfc3b;
#10;
address_ina = 162;
address_inb = 163;
data_ina = 16'h303;
data_inb = 16'hff37;
#10;
address_ina = 164;
address_inb = 165;
data_ina = 16'h50;
data_inb = 16'hf9b8;
#10;
address_ina = 166;
address_inb = 167;
data_ina = 16'h633;
data_inb = 16'hfe11;
#10;
address_ina = 168;
address_inb = 169;
data_ina = 16'hff1e;
data_inb = 16'hfc48;
#10;
address_ina = 170;
address_inb = 171;
data_ina = 16'hfa1c;
data_inb = 16'hf9c6;
#10;
address_ina = 172;
address_inb = 173;
data_ina = 16'h5f3;
data_inb = 16'h666;
#10;
address_ina = 174;
address_inb = 175;
data_ina = 16'h15e;
data_inb = 16'h1a5;
#10;
address_ina = 176;
address_inb = 177;
data_ina = 16'hfed5;
data_inb = 16'hfbfd;
#10;
address_ina = 178;
address_inb = 179;
data_ina = 16'h5fd;
data_inb = 16'h507;
#10;
address_ina = 180;
address_inb = 181;
data_ina = 16'hfa83;
data_inb = 16'hff18;
#10;
address_ina = 182;
address_inb = 183;
data_ina = 16'h9;
data_inb = 16'hfcba;
#10;
address_ina = 184;
address_inb = 185;
data_ina = 16'h290;
data_inb = 16'hfce8;
#10;
address_ina = 186;
address_inb = 187;
data_ina = 16'hfb2f;
data_inb = 16'hfdac;
#10;
address_ina = 188;
address_inb = 189;
data_ina = 16'hfd68;
data_inb = 16'hfea9;
#10;
address_ina = 190;
address_inb = 191;
data_ina = 16'h3c7;
data_inb = 16'h45a;
#10;
address_ina = 192;
address_inb = 193;
data_ina = 16'hfc4d;
data_inb = 16'hfa8a;
#10;
address_ina = 194;
address_inb = 195;
data_ina = 16'h2ad;
data_inb = 16'hfcfe;
#10;
address_ina = 196;
address_inb = 197;
data_ina = 16'h33f;
data_inb = 16'hfb04;
#10;
address_ina = 198;
address_inb = 199;
data_ina = 16'hfeaf;
data_inb = 16'hfa3d;
#10;
address_ina = 200;
address_inb = 201;
data_ina = 16'h601;
data_inb = 16'h3cb;
#10;
address_ina = 202;
address_inb = 203;
data_ina = 16'h40c;
data_inb = 16'h67;
#10;
address_ina = 204;
address_inb = 205;
data_ina = 16'hfbf0;
data_inb = 16'hb7;
#10;
address_ina = 206;
address_inb = 207;
data_ina = 16'hff8b;
data_inb = 16'hfc6b;
#10;
address_ina = 208;
address_inb = 209;
data_ina = 16'h396;
data_inb = 16'h363;
#10;
address_ina = 210;
address_inb = 211;
data_ina = 16'hfc53;
data_inb = 16'hff01;
#10;
address_ina = 212;
address_inb = 213;
data_ina = 16'hfee7;
data_inb = 16'h190;
#10;
address_ina = 214;
address_inb = 215;
data_ina = 16'h492;
data_inb = 16'h8b;
#10;
address_ina = 216;
address_inb = 217;
data_ina = 16'hff9b;
data_inb = 16'hfdfd;
#10;
address_ina = 218;
address_inb = 219;
data_ina = 16'he7;
data_inb = 16'h675;
#10;
address_ina = 220;
address_inb = 221;
data_ina = 16'h24a;
data_inb = 16'h26a;
#10;
address_ina = 222;
address_inb = 223;
data_ina = 16'h4fd;
data_inb = 16'h284;
#10;
address_ina = 224;
address_inb = 225;
data_ina = 16'hfab6;
data_inb = 16'hfc5f;
#10;
address_ina = 226;
address_inb = 227;
data_ina = 16'hfc6b;
data_inb = 16'h4fe;
#10;
address_ina = 228;
address_inb = 229;
data_ina = 16'h295;
data_inb = 16'hfe96;
#10;
address_ina = 230;
address_inb = 231;
data_ina = 16'hfb96;
data_inb = 16'hfeac;
#10;
address_ina = 232;
address_inb = 233;
data_ina = 16'hf4;
data_inb = 16'h9d;
#10;
address_ina = 234;
address_inb = 235;
data_ina = 16'hfb27;
data_inb = 16'hfd89;
#10;
address_ina = 236;
address_inb = 237;
data_ina = 16'h1b3;
data_inb = 16'hd9;
#10;
address_ina = 238;
address_inb = 239;
data_ina = 16'h171;
data_inb = 16'hfb45;
#10;
address_ina = 240;
address_inb = 241;
data_ina = 16'hfffb;
data_inb = 16'hf985;
#10;
address_ina = 242;
address_inb = 243;
data_ina = 16'h400;
data_inb = 16'hfc81;
#10;
address_ina = 244;
address_inb = 245;
data_ina = 16'hfd6f;
data_inb = 16'h39a;
#10;
address_ina = 246;
address_inb = 247;
data_ina = 16'h4dd;
data_inb = 16'hfb0b;
#10;
address_ina = 248;
address_inb = 249;
data_ina = 16'hfaad;
data_inb = 16'hf9ab;
#10;
address_ina = 250;
address_inb = 251;
data_ina = 16'h599;
data_inb = 16'h44f;
#10;
address_ina = 252;
address_inb = 253;
data_ina = 16'h4dc;
data_inb = 16'hfc75;
#10;
address_ina = 254;
address_inb = 255;
data_ina = 16'h59c;
data_inb = 16'h1ec;
#10;
        wait(init_done);
        #30
        we = 0;
        // Start processing
         
		  #38000

        start = 0;



//        wait (wr_req);
//		  wait (!wr_req);
//		   rd_req = 1;
		  wait(done);
		  #20000
rd_req = 1;
        #70 
		  start = 1;
		 #80 
wait(rd_empty)
rd_req = 0;

$display("Finished the NTT test Number %d",test_num);
////Begin test number #66//////////////
rst = 1;

//#1000
start = 1;
mode = 1; //NTT 0 // INTT 1

// Reset for a few clock cycles

#1000

rst = 0;
test_num = test_num + 1;
#1000
we = 1;
address_ina = 0;
address_inb = 1;
data_ina = 16'hfd7b;
data_inb = 16'hfd91;
#10;
address_ina = 2;
address_inb = 3;
data_ina = 16'h5da;
data_inb = 16'h24c;
#10;
address_ina = 4;
address_inb = 5;
data_ina = 16'h59b;
data_inb = 16'h64a;
#10;
address_ina = 6;
address_inb = 7;
data_ina = 16'h594;
data_inb = 16'hfad7;
#10;
address_ina = 8;
address_inb = 9;
data_ina = 16'hf993;
data_inb = 16'h2b2;
#10;
address_ina = 10;
address_inb = 11;
data_ina = 16'ha;
data_inb = 16'hffcc;
#10;
address_ina = 12;
address_inb = 13;
data_ina = 16'hfeb7;
data_inb = 16'hf9d8;
#10;
address_ina = 14;
address_inb = 15;
data_ina = 16'h3ae;
data_inb = 16'hfd50;
#10;
address_ina = 16;
address_inb = 17;
data_ina = 16'h550;
data_inb = 16'hf9a2;
#10;
address_ina = 18;
address_inb = 19;
data_ina = 16'hfceb;
data_inb = 16'h567;
#10;
address_ina = 20;
address_inb = 21;
data_ina = 16'h121;
data_inb = 16'h182;
#10;
address_ina = 22;
address_inb = 23;
data_ina = 16'h65f;
data_inb = 16'h4bf;
#10;
address_ina = 24;
address_inb = 25;
data_ina = 16'h135;
data_inb = 16'hde;
#10;
address_ina = 26;
address_inb = 27;
data_ina = 16'hfd7b;
data_inb = 16'h272;
#10;
address_ina = 28;
address_inb = 29;
data_ina = 16'h4ae;
data_inb = 16'h2ff;
#10;
address_ina = 30;
address_inb = 31;
data_ina = 16'hfa78;
data_inb = 16'h329;
#10;
address_ina = 32;
address_inb = 33;
data_ina = 16'hfc08;
data_inb = 16'h2ad;
#10;
address_ina = 34;
address_inb = 35;
data_ina = 16'hfa77;
data_inb = 16'hffbb;
#10;
address_ina = 36;
address_inb = 37;
data_ina = 16'hfe09;
data_inb = 16'hfb4d;
#10;
address_ina = 38;
address_inb = 39;
data_ina = 16'h502;
data_inb = 16'h1d6;
#10;
address_ina = 40;
address_inb = 41;
data_ina = 16'hfe48;
data_inb = 16'hffbd;
#10;
address_ina = 42;
address_inb = 43;
data_ina = 16'hfae6;
data_inb = 16'hfbbc;
#10;
address_ina = 44;
address_inb = 45;
data_ina = 16'h2ac;
data_inb = 16'h48c;
#10;
address_ina = 46;
address_inb = 47;
data_ina = 16'h3f6;
data_inb = 16'hfb3d;
#10;
address_ina = 48;
address_inb = 49;
data_ina = 16'hfbb3;
data_inb = 16'hfd24;
#10;
address_ina = 50;
address_inb = 51;
data_ina = 16'hfd44;
data_inb = 16'h318;
#10;
address_ina = 52;
address_inb = 53;
data_ina = 16'h44;
data_inb = 16'h660;
#10;
address_ina = 54;
address_inb = 55;
data_ina = 16'hfe6e;
data_inb = 16'hfe97;
#10;
address_ina = 56;
address_inb = 57;
data_ina = 16'hfe99;
data_inb = 16'h37c;
#10;
address_ina = 58;
address_inb = 59;
data_ina = 16'hfca0;
data_inb = 16'h593;
#10;
address_ina = 60;
address_inb = 61;
data_ina = 16'h283;
data_inb = 16'h1a5;
#10;
address_ina = 62;
address_inb = 63;
data_ina = 16'h80;
data_inb = 16'hfce0;
#10;
address_ina = 64;
address_inb = 65;
data_ina = 16'hf99e;
data_inb = 16'h53b;
#10;
address_ina = 66;
address_inb = 67;
data_ina = 16'h62d;
data_inb = 16'hff6f;
#10;
address_ina = 68;
address_inb = 69;
data_ina = 16'h408;
data_inb = 16'hff96;
#10;
address_ina = 70;
address_inb = 71;
data_ina = 16'h13f;
data_inb = 16'hfa23;
#10;
address_ina = 72;
address_inb = 73;
data_ina = 16'h1d6;
data_inb = 16'h53e;
#10;
address_ina = 74;
address_inb = 75;
data_ina = 16'hfd73;
data_inb = 16'hf989;
#10;
address_ina = 76;
address_inb = 77;
data_ina = 16'hfc97;
data_inb = 16'h241;
#10;
address_ina = 78;
address_inb = 79;
data_ina = 16'h375;
data_inb = 16'hff3e;
#10;
address_ina = 80;
address_inb = 81;
data_ina = 16'h574;
data_inb = 16'hfbd5;
#10;
address_ina = 82;
address_inb = 83;
data_ina = 16'h184;
data_inb = 16'h58f;
#10;
address_ina = 84;
address_inb = 85;
data_ina = 16'he7;
data_inb = 16'hfae1;
#10;
address_ina = 86;
address_inb = 87;
data_ina = 16'h137;
data_inb = 16'h1ad;
#10;
address_ina = 88;
address_inb = 89;
data_ina = 16'hfa13;
data_inb = 16'h15;
#10;
address_ina = 90;
address_inb = 91;
data_ina = 16'h48;
data_inb = 16'hfde1;
#10;
address_ina = 92;
address_inb = 93;
data_ina = 16'h203;
data_inb = 16'h3c7;
#10;
address_ina = 94;
address_inb = 95;
data_ina = 16'h433;
data_inb = 16'hfdff;
#10;
address_ina = 96;
address_inb = 97;
data_ina = 16'h545;
data_inb = 16'hfc5b;
#10;
address_ina = 98;
address_inb = 99;
data_ina = 16'hff9c;
data_inb = 16'h146;
#10;
address_ina = 100;
address_inb = 101;
data_ina = 16'h3a5;
data_inb = 16'hfdea;
#10;
address_ina = 102;
address_inb = 103;
data_ina = 16'h254;
data_inb = 16'h2a6;
#10;
address_ina = 104;
address_inb = 105;
data_ina = 16'hfba4;
data_inb = 16'h40;
#10;
address_ina = 106;
address_inb = 107;
data_ina = 16'h12;
data_inb = 16'h3a9;
#10;
address_ina = 108;
address_inb = 109;
data_ina = 16'h5fd;
data_inb = 16'h2e;
#10;
address_ina = 110;
address_inb = 111;
data_ina = 16'hfd58;
data_inb = 16'hffa6;
#10;
address_ina = 112;
address_inb = 113;
data_ina = 16'h424;
data_inb = 16'hfc4c;
#10;
address_ina = 114;
address_inb = 115;
data_ina = 16'h305;
data_inb = 16'h2bb;
#10;
address_ina = 116;
address_inb = 117;
data_ina = 16'h30a;
data_inb = 16'hfc37;
#10;
address_ina = 118;
address_inb = 119;
data_ina = 16'h13e;
data_inb = 16'h13;
#10;
address_ina = 120;
address_inb = 121;
data_ina = 16'h5e;
data_inb = 16'hfcc5;
#10;
address_ina = 122;
address_inb = 123;
data_ina = 16'h1c2;
data_inb = 16'hfd53;
#10;
address_ina = 124;
address_inb = 125;
data_ina = 16'hfb7e;
data_inb = 16'hfc93;
#10;
address_ina = 126;
address_inb = 127;
data_ina = 16'h5dc;
data_inb = 16'hfe89;
#10;
address_ina = 128;
address_inb = 129;
data_ina = 16'h2a1;
data_inb = 16'h153;
#10;
address_ina = 130;
address_inb = 131;
data_ina = 16'hfb2e;
data_inb = 16'hfb06;
#10;
address_ina = 132;
address_inb = 133;
data_ina = 16'hfe4e;
data_inb = 16'h252;
#10;
address_ina = 134;
address_inb = 135;
data_ina = 16'h55f;
data_inb = 16'h5ae;
#10;
address_ina = 136;
address_inb = 137;
data_ina = 16'h258;
data_inb = 16'hff8b;
#10;
address_ina = 138;
address_inb = 139;
data_ina = 16'h152;
data_inb = 16'hfe9d;
#10;
address_ina = 140;
address_inb = 141;
data_ina = 16'hfab3;
data_inb = 16'hfdb7;
#10;
address_ina = 142;
address_inb = 143;
data_ina = 16'h3b;
data_inb = 16'hfb3f;
#10;
address_ina = 144;
address_inb = 145;
data_ina = 16'h27b;
data_inb = 16'h432;
#10;
address_ina = 146;
address_inb = 147;
data_ina = 16'hfd47;
data_inb = 16'hfb61;
#10;
address_ina = 148;
address_inb = 149;
data_ina = 16'hfc9d;
data_inb = 16'h12a;
#10;
address_ina = 150;
address_inb = 151;
data_ina = 16'h5ec;
data_inb = 16'h313;
#10;
address_ina = 152;
address_inb = 153;
data_ina = 16'h639;
data_inb = 16'hfc0d;
#10;
address_ina = 154;
address_inb = 155;
data_ina = 16'hfcf5;
data_inb = 16'hfa88;
#10;
address_ina = 156;
address_inb = 157;
data_ina = 16'h340;
data_inb = 16'hfa63;
#10;
address_ina = 158;
address_inb = 159;
data_ina = 16'h596;
data_inb = 16'h5d9;
#10;
address_ina = 160;
address_inb = 161;
data_ina = 16'hfaa0;
data_inb = 16'hfb32;
#10;
address_ina = 162;
address_inb = 163;
data_ina = 16'h2ef;
data_inb = 16'hfece;
#10;
address_ina = 164;
address_inb = 165;
data_ina = 16'h23b;
data_inb = 16'h35a;
#10;
address_ina = 166;
address_inb = 167;
data_ina = 16'hfbfa;
data_inb = 16'h84;
#10;
address_ina = 168;
address_inb = 169;
data_ina = 16'h224;
data_inb = 16'h4bc;
#10;
address_ina = 170;
address_inb = 171;
data_ina = 16'h3a3;
data_inb = 16'hfe72;
#10;
address_ina = 172;
address_inb = 173;
data_ina = 16'hf9c5;
data_inb = 16'h50b;
#10;
address_ina = 174;
address_inb = 175;
data_ina = 16'h2cf;
data_inb = 16'hfaed;
#10;
address_ina = 176;
address_inb = 177;
data_ina = 16'h3e0;
data_inb = 16'h3a0;
#10;
address_ina = 178;
address_inb = 179;
data_ina = 16'h3cc;
data_inb = 16'hff3b;
#10;
address_ina = 180;
address_inb = 181;
data_ina = 16'h42c;
data_inb = 16'hfc14;
#10;
address_ina = 182;
address_inb = 183;
data_ina = 16'h5c1;
data_inb = 16'h524;
#10;
address_ina = 184;
address_inb = 185;
data_ina = 16'h36d;
data_inb = 16'h422;
#10;
address_ina = 186;
address_inb = 187;
data_ina = 16'h21a;
data_inb = 16'hfef0;
#10;
address_ina = 188;
address_inb = 189;
data_ina = 16'hfad8;
data_inb = 16'h219;
#10;
address_ina = 190;
address_inb = 191;
data_ina = 16'hfcb0;
data_inb = 16'h82;
#10;
address_ina = 192;
address_inb = 193;
data_ina = 16'hfd8e;
data_inb = 16'h2fd;
#10;
address_ina = 194;
address_inb = 195;
data_ina = 16'h104;
data_inb = 16'h120;
#10;
address_ina = 196;
address_inb = 197;
data_ina = 16'hfeab;
data_inb = 16'h49a;
#10;
address_ina = 198;
address_inb = 199;
data_ina = 16'h129;
data_inb = 16'hfa9b;
#10;
address_ina = 200;
address_inb = 201;
data_ina = 16'h1a8;
data_inb = 16'hfbed;
#10;
address_ina = 202;
address_inb = 203;
data_ina = 16'hfe31;
data_inb = 16'hfd60;
#10;
address_ina = 204;
address_inb = 205;
data_ina = 16'h333;
data_inb = 16'h538;
#10;
address_ina = 206;
address_inb = 207;
data_ina = 16'hfa45;
data_inb = 16'hfb91;
#10;
address_ina = 208;
address_inb = 209;
data_ina = 16'hff62;
data_inb = 16'hfbfe;
#10;
address_ina = 210;
address_inb = 211;
data_ina = 16'h344;
data_inb = 16'hfef2;
#10;
address_ina = 212;
address_inb = 213;
data_ina = 16'h61b;
data_inb = 16'hfec2;
#10;
address_ina = 214;
address_inb = 215;
data_ina = 16'hff97;
data_inb = 16'hfd80;
#10;
address_ina = 216;
address_inb = 217;
data_ina = 16'hff10;
data_inb = 16'hfb87;
#10;
address_ina = 218;
address_inb = 219;
data_ina = 16'hff3f;
data_inb = 16'h3e8;
#10;
address_ina = 220;
address_inb = 221;
data_ina = 16'hfdd9;
data_inb = 16'hfeec;
#10;
address_ina = 222;
address_inb = 223;
data_ina = 16'hfcf7;
data_inb = 16'hffbf;
#10;
address_ina = 224;
address_inb = 225;
data_ina = 16'hfc79;
data_inb = 16'h10c;
#10;
address_ina = 226;
address_inb = 227;
data_ina = 16'h5d1;
data_inb = 16'h26b;
#10;
address_ina = 228;
address_inb = 229;
data_ina = 16'h3be;
data_inb = 16'h4cb;
#10;
address_ina = 230;
address_inb = 231;
data_ina = 16'h119;
data_inb = 16'h436;
#10;
address_ina = 232;
address_inb = 233;
data_ina = 16'hfb68;
data_inb = 16'h4f8;
#10;
address_ina = 234;
address_inb = 235;
data_ina = 16'hfbf0;
data_inb = 16'h531;
#10;
address_ina = 236;
address_inb = 237;
data_ina = 16'hfd60;
data_inb = 16'hfccb;
#10;
address_ina = 238;
address_inb = 239;
data_ina = 16'h182;
data_inb = 16'h653;
#10;
address_ina = 240;
address_inb = 241;
data_ina = 16'hfe06;
data_inb = 16'hfe8b;
#10;
address_ina = 242;
address_inb = 243;
data_ina = 16'h393;
data_inb = 16'hfdaf;
#10;
address_ina = 244;
address_inb = 245;
data_ina = 16'hff9a;
data_inb = 16'hff80;
#10;
address_ina = 246;
address_inb = 247;
data_ina = 16'hfe05;
data_inb = 16'h133;
#10;
address_ina = 248;
address_inb = 249;
data_ina = 16'h323;
data_inb = 16'hfb1f;
#10;
address_ina = 250;
address_inb = 251;
data_ina = 16'hf9e8;
data_inb = 16'h2f7;
#10;
address_ina = 252;
address_inb = 253;
data_ina = 16'hfab4;
data_inb = 16'h39e;
#10;
address_ina = 254;
address_inb = 255;
data_ina = 16'hfeb3;
data_inb = 16'h268;
#10;
        wait(init_done);
        #30
        we = 0;
        // Start processing
         
		  #38000

        start = 0;



//        wait (wr_req);
//		  wait (!wr_req);
//		   rd_req = 1;
		  wait(done);
		  #20000
rd_req = 1;
        #70 
		  start = 1;
		 #80 
wait(rd_empty)
rd_req = 0;

$display("Finished the NTT test Number %d",test_num);
////Begin test number #67//////////////
rst = 1;

//#1000
start = 1;
mode = 1; //NTT 0 // INTT 1

// Reset for a few clock cycles

#1000

rst = 0;
test_num = test_num + 1;
#1000
we = 1;
address_ina = 0;
address_inb = 1;
data_ina = 16'hff7d;
data_inb = 16'h2c8;
#10;
address_ina = 2;
address_inb = 3;
data_ina = 16'hfcf9;
data_inb = 16'hfaa6;
#10;
address_ina = 4;
address_inb = 5;
data_ina = 16'h58;
data_inb = 16'h43c;
#10;
address_ina = 6;
address_inb = 7;
data_ina = 16'h23e;
data_inb = 16'hfaa2;
#10;
address_ina = 8;
address_inb = 9;
data_ina = 16'hff48;
data_inb = 16'h1dc;
#10;
address_ina = 10;
address_inb = 11;
data_ina = 16'h5d3;
data_inb = 16'hfdc0;
#10;
address_ina = 12;
address_inb = 13;
data_ina = 16'hfce1;
data_inb = 16'h5e1;
#10;
address_ina = 14;
address_inb = 15;
data_ina = 16'h66e;
data_inb = 16'h3c3;
#10;
address_ina = 16;
address_inb = 17;
data_ina = 16'hfe10;
data_inb = 16'hfb44;
#10;
address_ina = 18;
address_inb = 19;
data_ina = 16'h278;
data_inb = 16'hfbac;
#10;
address_ina = 20;
address_inb = 21;
data_ina = 16'hfe40;
data_inb = 16'h442;
#10;
address_ina = 22;
address_inb = 23;
data_ina = 16'hff62;
data_inb = 16'hfda7;
#10;
address_ina = 24;
address_inb = 25;
data_ina = 16'h4e;
data_inb = 16'heb;
#10;
address_ina = 26;
address_inb = 27;
data_ina = 16'h35e;
data_inb = 16'h26e;
#10;
address_ina = 28;
address_inb = 29;
data_ina = 16'hfc2c;
data_inb = 16'h4bb;
#10;
address_ina = 30;
address_inb = 31;
data_ina = 16'h28;
data_inb = 16'hfb60;
#10;
address_ina = 32;
address_inb = 33;
data_ina = 16'hfb1d;
data_inb = 16'h41d;
#10;
address_ina = 34;
address_inb = 35;
data_ina = 16'hfc79;
data_inb = 16'h426;
#10;
address_ina = 36;
address_inb = 37;
data_ina = 16'hfb75;
data_inb = 16'h193;
#10;
address_ina = 38;
address_inb = 39;
data_ina = 16'hfcc1;
data_inb = 16'hfeb0;
#10;
address_ina = 40;
address_inb = 41;
data_ina = 16'h164;
data_inb = 16'h5fa;
#10;
address_ina = 42;
address_inb = 43;
data_ina = 16'h37;
data_inb = 16'hfd86;
#10;
address_ina = 44;
address_inb = 45;
data_ina = 16'hfe9e;
data_inb = 16'hfee9;
#10;
address_ina = 46;
address_inb = 47;
data_ina = 16'h3f1;
data_inb = 16'h623;
#10;
address_ina = 48;
address_inb = 49;
data_ina = 16'hfd3e;
data_inb = 16'hfde8;
#10;
address_ina = 50;
address_inb = 51;
data_ina = 16'hfc89;
data_inb = 16'h4d8;
#10;
address_ina = 52;
address_inb = 53;
data_ina = 16'hfcbd;
data_inb = 16'hfb3b;
#10;
address_ina = 54;
address_inb = 55;
data_ina = 16'h609;
data_inb = 16'hfd3d;
#10;
address_ina = 56;
address_inb = 57;
data_ina = 16'h134;
data_inb = 16'hffe9;
#10;
address_ina = 58;
address_inb = 59;
data_ina = 16'hff64;
data_inb = 16'h29f;
#10;
address_ina = 60;
address_inb = 61;
data_ina = 16'h1ec;
data_inb = 16'h5c5;
#10;
address_ina = 62;
address_inb = 63;
data_ina = 16'h4fd;
data_inb = 16'h187;
#10;
address_ina = 64;
address_inb = 65;
data_ina = 16'hf9e4;
data_inb = 16'h303;
#10;
address_ina = 66;
address_inb = 67;
data_ina = 16'h40f;
data_inb = 16'h13d;
#10;
address_ina = 68;
address_inb = 69;
data_ina = 16'hff29;
data_inb = 16'h2c9;
#10;
address_ina = 70;
address_inb = 71;
data_ina = 16'hfec9;
data_inb = 16'hfec0;
#10;
address_ina = 72;
address_inb = 73;
data_ina = 16'hfde5;
data_inb = 16'hfdaa;
#10;
address_ina = 74;
address_inb = 75;
data_ina = 16'h258;
data_inb = 16'hfc14;
#10;
address_ina = 76;
address_inb = 77;
data_ina = 16'h434;
data_inb = 16'hf9f7;
#10;
address_ina = 78;
address_inb = 79;
data_ina = 16'hff65;
data_inb = 16'hff04;
#10;
address_ina = 80;
address_inb = 81;
data_ina = 16'hfdcb;
data_inb = 16'hf9b4;
#10;
address_ina = 82;
address_inb = 83;
data_ina = 16'h163;
data_inb = 16'hfcf2;
#10;
address_ina = 84;
address_inb = 85;
data_ina = 16'h602;
data_inb = 16'hfd73;
#10;
address_ina = 86;
address_inb = 87;
data_ina = 16'hfa17;
data_inb = 16'h384;
#10;
address_ina = 88;
address_inb = 89;
data_ina = 16'h2c6;
data_inb = 16'h323;
#10;
address_ina = 90;
address_inb = 91;
data_ina = 16'h3d;
data_inb = 16'hfeb5;
#10;
address_ina = 92;
address_inb = 93;
data_ina = 16'h331;
data_inb = 16'h367;
#10;
address_ina = 94;
address_inb = 95;
data_ina = 16'hfaa2;
data_inb = 16'hfcd6;
#10;
address_ina = 96;
address_inb = 97;
data_ina = 16'hfad8;
data_inb = 16'h3b2;
#10;
address_ina = 98;
address_inb = 99;
data_ina = 16'h1a9;
data_inb = 16'h568;
#10;
address_ina = 100;
address_inb = 101;
data_ina = 16'hfdb5;
data_inb = 16'hfa87;
#10;
address_ina = 102;
address_inb = 103;
data_ina = 16'h46;
data_inb = 16'hfc3a;
#10;
address_ina = 104;
address_inb = 105;
data_ina = 16'h1ec;
data_inb = 16'h18a;
#10;
address_ina = 106;
address_inb = 107;
data_ina = 16'h436;
data_inb = 16'hf9b2;
#10;
address_ina = 108;
address_inb = 109;
data_ina = 16'hff99;
data_inb = 16'h2d2;
#10;
address_ina = 110;
address_inb = 111;
data_ina = 16'hffee;
data_inb = 16'h30f;
#10;
address_ina = 112;
address_inb = 113;
data_ina = 16'h1f1;
data_inb = 16'hfda7;
#10;
address_ina = 114;
address_inb = 115;
data_ina = 16'h609;
data_inb = 16'h4f9;
#10;
address_ina = 116;
address_inb = 117;
data_ina = 16'hfa84;
data_inb = 16'hff22;
#10;
address_ina = 118;
address_inb = 119;
data_ina = 16'hfd67;
data_inb = 16'h319;
#10;
address_ina = 120;
address_inb = 121;
data_ina = 16'hfb17;
data_inb = 16'hfa43;
#10;
address_ina = 122;
address_inb = 123;
data_ina = 16'h4e0;
data_inb = 16'h2e7;
#10;
address_ina = 124;
address_inb = 125;
data_ina = 16'hfb5d;
data_inb = 16'hfe49;
#10;
address_ina = 126;
address_inb = 127;
data_ina = 16'h384;
data_inb = 16'h395;
#10;
address_ina = 128;
address_inb = 129;
data_ina = 16'h160;
data_inb = 16'hffff;
#10;
address_ina = 130;
address_inb = 131;
data_ina = 16'h390;
data_inb = 16'h2f1;
#10;
address_ina = 132;
address_inb = 133;
data_ina = 16'h4aa;
data_inb = 16'hf9c6;
#10;
address_ina = 134;
address_inb = 135;
data_ina = 16'hfe46;
data_inb = 16'hfefb;
#10;
address_ina = 136;
address_inb = 137;
data_ina = 16'hfd0e;
data_inb = 16'h217;
#10;
address_ina = 138;
address_inb = 139;
data_ina = 16'hfc8f;
data_inb = 16'h321;
#10;
address_ina = 140;
address_inb = 141;
data_ina = 16'h467;
data_inb = 16'hfd70;
#10;
address_ina = 142;
address_inb = 143;
data_ina = 16'h1db;
data_inb = 16'h628;
#10;
address_ina = 144;
address_inb = 145;
data_ina = 16'h5ba;
data_inb = 16'h421;
#10;
address_ina = 146;
address_inb = 147;
data_ina = 16'hfc1f;
data_inb = 16'hffeb;
#10;
address_ina = 148;
address_inb = 149;
data_ina = 16'hfd0e;
data_inb = 16'h455;
#10;
address_ina = 150;
address_inb = 151;
data_ina = 16'hfa41;
data_inb = 16'h182;
#10;
address_ina = 152;
address_inb = 153;
data_ina = 16'hfd94;
data_inb = 16'hfc0f;
#10;
address_ina = 154;
address_inb = 155;
data_ina = 16'hfe8e;
data_inb = 16'hfb66;
#10;
address_ina = 156;
address_inb = 157;
data_ina = 16'h4d7;
data_inb = 16'h27f;
#10;
address_ina = 158;
address_inb = 159;
data_ina = 16'h17f;
data_inb = 16'hab;
#10;
address_ina = 160;
address_inb = 161;
data_ina = 16'h36a;
data_inb = 16'hea;
#10;
address_ina = 162;
address_inb = 163;
data_ina = 16'ha1;
data_inb = 16'h467;
#10;
address_ina = 164;
address_inb = 165;
data_ina = 16'h2ed;
data_inb = 16'h53a;
#10;
address_ina = 166;
address_inb = 167;
data_ina = 16'h68;
data_inb = 16'hfc9c;
#10;
address_ina = 168;
address_inb = 169;
data_ina = 16'hfc4d;
data_inb = 16'h578;
#10;
address_ina = 170;
address_inb = 171;
data_ina = 16'h34f;
data_inb = 16'h5a4;
#10;
address_ina = 172;
address_inb = 173;
data_ina = 16'hab;
data_inb = 16'hfc2e;
#10;
address_ina = 174;
address_inb = 175;
data_ina = 16'hfc13;
data_inb = 16'hfec2;
#10;
address_ina = 176;
address_inb = 177;
data_ina = 16'h1af;
data_inb = 16'hfa73;
#10;
address_ina = 178;
address_inb = 179;
data_ina = 16'hfc44;
data_inb = 16'hfb6c;
#10;
address_ina = 180;
address_inb = 181;
data_ina = 16'h541;
data_inb = 16'hfe84;
#10;
address_ina = 182;
address_inb = 183;
data_ina = 16'h359;
data_inb = 16'h24c;
#10;
address_ina = 184;
address_inb = 185;
data_ina = 16'hfe2b;
data_inb = 16'h2b;
#10;
address_ina = 186;
address_inb = 187;
data_ina = 16'hfcf9;
data_inb = 16'h4f5;
#10;
address_ina = 188;
address_inb = 189;
data_ina = 16'h66d;
data_inb = 16'hff69;
#10;
address_ina = 190;
address_inb = 191;
data_ina = 16'hfd47;
data_inb = 16'h3f;
#10;
address_ina = 192;
address_inb = 193;
data_ina = 16'h18a;
data_inb = 16'hfa8d;
#10;
address_ina = 194;
address_inb = 195;
data_ina = 16'h4cd;
data_inb = 16'hf9;
#10;
address_ina = 196;
address_inb = 197;
data_ina = 16'h331;
data_inb = 16'hfb91;
#10;
address_ina = 198;
address_inb = 199;
data_ina = 16'h38a;
data_inb = 16'h362;
#10;
address_ina = 200;
address_inb = 201;
data_ina = 16'h18d;
data_inb = 16'h680;
#10;
address_ina = 202;
address_inb = 203;
data_ina = 16'hfb3f;
data_inb = 16'hfb64;
#10;
address_ina = 204;
address_inb = 205;
data_ina = 16'hfe83;
data_inb = 16'h42b;
#10;
address_ina = 206;
address_inb = 207;
data_ina = 16'hfa1b;
data_inb = 16'h59c;
#10;
address_ina = 208;
address_inb = 209;
data_ina = 16'hffe5;
data_inb = 16'h586;
#10;
address_ina = 210;
address_inb = 211;
data_ina = 16'h374;
data_inb = 16'hd6;
#10;
address_ina = 212;
address_inb = 213;
data_ina = 16'h74;
data_inb = 16'hfba6;
#10;
address_ina = 214;
address_inb = 215;
data_ina = 16'h4c3;
data_inb = 16'h34f;
#10;
address_ina = 216;
address_inb = 217;
data_ina = 16'h41c;
data_inb = 16'h2f;
#10;
address_ina = 218;
address_inb = 219;
data_ina = 16'h27e;
data_inb = 16'h3b5;
#10;
address_ina = 220;
address_inb = 221;
data_ina = 16'hff7e;
data_inb = 16'h61d;
#10;
address_ina = 222;
address_inb = 223;
data_ina = 16'hfd37;
data_inb = 16'hfed3;
#10;
address_ina = 224;
address_inb = 225;
data_ina = 16'h2fe;
data_inb = 16'hfb53;
#10;
address_ina = 226;
address_inb = 227;
data_ina = 16'hfe14;
data_inb = 16'hfb9c;
#10;
address_ina = 228;
address_inb = 229;
data_ina = 16'hfdeb;
data_inb = 16'h347;
#10;
address_ina = 230;
address_inb = 231;
data_ina = 16'hfcf9;
data_inb = 16'h575;
#10;
address_ina = 232;
address_inb = 233;
data_ina = 16'h549;
data_inb = 16'h163;
#10;
address_ina = 234;
address_inb = 235;
data_ina = 16'hfd8c;
data_inb = 16'hfae2;
#10;
address_ina = 236;
address_inb = 237;
data_ina = 16'h5cc;
data_inb = 16'h2e;
#10;
address_ina = 238;
address_inb = 239;
data_ina = 16'h397;
data_inb = 16'hfab9;
#10;
address_ina = 240;
address_inb = 241;
data_ina = 16'h1bb;
data_inb = 16'h24;
#10;
address_ina = 242;
address_inb = 243;
data_ina = 16'hff1d;
data_inb = 16'hf9a0;
#10;
address_ina = 244;
address_inb = 245;
data_ina = 16'h651;
data_inb = 16'hfb13;
#10;
address_ina = 246;
address_inb = 247;
data_ina = 16'h5f8;
data_inb = 16'hfb03;
#10;
address_ina = 248;
address_inb = 249;
data_ina = 16'hfd74;
data_inb = 16'h142;
#10;
address_ina = 250;
address_inb = 251;
data_ina = 16'h566;
data_inb = 16'hfa6a;
#10;
address_ina = 252;
address_inb = 253;
data_ina = 16'hff97;
data_inb = 16'hfd24;
#10;
address_ina = 254;
address_inb = 255;
data_ina = 16'h2a0;
data_inb = 16'h5ef;
#10;
        wait(init_done);
        #30
        we = 0;
        // Start processing
         
		  #38000

        start = 0;



//        wait (wr_req);
//		  wait (!wr_req);
//		   rd_req = 1;
		  wait(done);
		  #20000
rd_req = 1;
        #70 
		  start = 1;
		 #80 
wait(rd_empty)
rd_req = 0;

$display("Finished the NTT test Number %d",test_num);
////Begin test number #68//////////////
rst = 1;

//#1000
start = 1;
mode = 0; //NTT 0 // INTT 1

// Reset for a few clock cycles

#1000

rst = 0;
test_num = test_num + 1;
#1000
we = 1;
address_ina = 0;
address_inb = 1;
data_ina = 16'hfffe;
data_inb = 16'h0;
#10;
address_ina = 2;
address_inb = 3;
data_ina = 16'h2;
data_inb = 16'hffff;
#10;
address_ina = 4;
address_inb = 5;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 6;
address_inb = 7;
data_ina = 16'h1;
data_inb = 16'hfffe;
#10;
address_ina = 8;
address_inb = 9;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 10;
address_inb = 11;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 12;
address_inb = 13;
data_ina = 16'hfffe;
data_inb = 16'h0;
#10;
address_ina = 14;
address_inb = 15;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 16;
address_inb = 17;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 18;
address_inb = 19;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 20;
address_inb = 21;
data_ina = 16'hfffe;
data_inb = 16'hffff;
#10;
address_ina = 22;
address_inb = 23;
data_ina = 16'hfffe;
data_inb = 16'hffff;
#10;
address_ina = 24;
address_inb = 25;
data_ina = 16'h2;
data_inb = 16'h1;
#10;
address_ina = 26;
address_inb = 27;
data_ina = 16'hffff;
data_inb = 16'hfffe;
#10;
address_ina = 28;
address_inb = 29;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 30;
address_inb = 31;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 32;
address_inb = 33;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 34;
address_inb = 35;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 36;
address_inb = 37;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 38;
address_inb = 39;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 40;
address_inb = 41;
data_ina = 16'h1;
data_inb = 16'h2;
#10;
address_ina = 42;
address_inb = 43;
data_ina = 16'hfffe;
data_inb = 16'h2;
#10;
address_ina = 44;
address_inb = 45;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 46;
address_inb = 47;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 48;
address_inb = 49;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 50;
address_inb = 51;
data_ina = 16'hfffe;
data_inb = 16'hffff;
#10;
address_ina = 52;
address_inb = 53;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 54;
address_inb = 55;
data_ina = 16'hfffe;
data_inb = 16'h1;
#10;
address_ina = 56;
address_inb = 57;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 58;
address_inb = 59;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 60;
address_inb = 61;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 62;
address_inb = 63;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 64;
address_inb = 65;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 66;
address_inb = 67;
data_ina = 16'h2;
data_inb = 16'hffff;
#10;
address_ina = 68;
address_inb = 69;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 70;
address_inb = 71;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 72;
address_inb = 73;
data_ina = 16'hfffe;
data_inb = 16'h0;
#10;
address_ina = 74;
address_inb = 75;
data_ina = 16'h2;
data_inb = 16'h0;
#10;
address_ina = 76;
address_inb = 77;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 78;
address_inb = 79;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 80;
address_inb = 81;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 82;
address_inb = 83;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 84;
address_inb = 85;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 86;
address_inb = 87;
data_ina = 16'hfffe;
data_inb = 16'h1;
#10;
address_ina = 88;
address_inb = 89;
data_ina = 16'hfffe;
data_inb = 16'h1;
#10;
address_ina = 90;
address_inb = 91;
data_ina = 16'h1;
data_inb = 16'hfffe;
#10;
address_ina = 92;
address_inb = 93;
data_ina = 16'h2;
data_inb = 16'h1;
#10;
address_ina = 94;
address_inb = 95;
data_ina = 16'h3;
data_inb = 16'h0;
#10;
address_ina = 96;
address_inb = 97;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 98;
address_inb = 99;
data_ina = 16'h2;
data_inb = 16'h1;
#10;
address_ina = 100;
address_inb = 101;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 102;
address_inb = 103;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 104;
address_inb = 105;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 106;
address_inb = 107;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 108;
address_inb = 109;
data_ina = 16'hffff;
data_inb = 16'h2;
#10;
address_ina = 110;
address_inb = 111;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 112;
address_inb = 113;
data_ina = 16'h0;
data_inb = 16'h3;
#10;
address_ina = 114;
address_inb = 115;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 116;
address_inb = 117;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 118;
address_inb = 119;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 120;
address_inb = 121;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 122;
address_inb = 123;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 124;
address_inb = 125;
data_ina = 16'h1;
data_inb = 16'h2;
#10;
address_ina = 126;
address_inb = 127;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 128;
address_inb = 129;
data_ina = 16'hffff;
data_inb = 16'h2;
#10;
address_ina = 130;
address_inb = 131;
data_ina = 16'hfffe;
data_inb = 16'h2;
#10;
address_ina = 132;
address_inb = 133;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 134;
address_inb = 135;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 136;
address_inb = 137;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 138;
address_inb = 139;
data_ina = 16'h0;
data_inb = 16'hfffe;
#10;
address_ina = 140;
address_inb = 141;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 142;
address_inb = 143;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 144;
address_inb = 145;
data_ina = 16'h1;
data_inb = 16'h2;
#10;
address_ina = 146;
address_inb = 147;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 148;
address_inb = 149;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 150;
address_inb = 151;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 152;
address_inb = 153;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 154;
address_inb = 155;
data_ina = 16'hfffe;
data_inb = 16'hffff;
#10;
address_ina = 156;
address_inb = 157;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 158;
address_inb = 159;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 160;
address_inb = 161;
data_ina = 16'hfffe;
data_inb = 16'hfffe;
#10;
address_ina = 162;
address_inb = 163;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 164;
address_inb = 165;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 166;
address_inb = 167;
data_ina = 16'h2;
data_inb = 16'hffff;
#10;
address_ina = 168;
address_inb = 169;
data_ina = 16'h0;
data_inb = 16'hfffe;
#10;
address_ina = 170;
address_inb = 171;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 172;
address_inb = 173;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 174;
address_inb = 175;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 176;
address_inb = 177;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 178;
address_inb = 179;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 180;
address_inb = 181;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 182;
address_inb = 183;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 184;
address_inb = 185;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 186;
address_inb = 187;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 188;
address_inb = 189;
data_ina = 16'hffff;
data_inb = 16'h2;
#10;
address_ina = 190;
address_inb = 191;
data_ina = 16'hfffe;
data_inb = 16'h1;
#10;
address_ina = 192;
address_inb = 193;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 194;
address_inb = 195;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 196;
address_inb = 197;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 198;
address_inb = 199;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 200;
address_inb = 201;
data_ina = 16'h2;
data_inb = 16'h1;
#10;
address_ina = 202;
address_inb = 203;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 204;
address_inb = 205;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 206;
address_inb = 207;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 208;
address_inb = 209;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 210;
address_inb = 211;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 212;
address_inb = 213;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 214;
address_inb = 215;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 216;
address_inb = 217;
data_ina = 16'hfffe;
data_inb = 16'h0;
#10;
address_ina = 218;
address_inb = 219;
data_ina = 16'h3;
data_inb = 16'h2;
#10;
address_ina = 220;
address_inb = 221;
data_ina = 16'h1;
data_inb = 16'hfffe;
#10;
address_ina = 222;
address_inb = 223;
data_ina = 16'h2;
data_inb = 16'hfffe;
#10;
address_ina = 224;
address_inb = 225;
data_ina = 16'h0;
data_inb = 16'hfffe;
#10;
address_ina = 226;
address_inb = 227;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 228;
address_inb = 229;
data_ina = 16'h0;
data_inb = 16'hfffe;
#10;
address_ina = 230;
address_inb = 231;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 232;
address_inb = 233;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 234;
address_inb = 235;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 236;
address_inb = 237;
data_ina = 16'h0;
data_inb = 16'hfffe;
#10;
address_ina = 238;
address_inb = 239;
data_ina = 16'h3;
data_inb = 16'h2;
#10;
address_ina = 240;
address_inb = 241;
data_ina = 16'h2;
data_inb = 16'hffff;
#10;
address_ina = 242;
address_inb = 243;
data_ina = 16'h1;
data_inb = 16'h2;
#10;
address_ina = 244;
address_inb = 245;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 246;
address_inb = 247;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 248;
address_inb = 249;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 250;
address_inb = 251;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 252;
address_inb = 253;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 254;
address_inb = 255;
data_ina = 16'h0;
data_inb = 16'hfffd;
#10;
        wait(init_done);
        #30
        we = 0;
        // Start processing
         
		  #38000

        start = 0;



//        wait (wr_req);
//		  wait (!wr_req);
//		   rd_req = 1;
		  wait(done);
		  #20000
rd_req = 1;
        #70 
		  start = 1;
		 #80 
wait(rd_empty)
rd_req = 0;

$display("Finished the NTT test Number %d",test_num);
////Begin test number #69//////////////
rst = 1;

//#1000
start = 1;
mode = 0; //NTT 0 // INTT 1

// Reset for a few clock cycles

#1000

rst = 0;
test_num = test_num + 1;
#1000
we = 1;
address_ina = 0;
address_inb = 1;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 2;
address_inb = 3;
data_ina = 16'hffff;
data_inb = 16'h2;
#10;
address_ina = 4;
address_inb = 5;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 6;
address_inb = 7;
data_ina = 16'hfffe;
data_inb = 16'h0;
#10;
address_ina = 8;
address_inb = 9;
data_ina = 16'h3;
data_inb = 16'h1;
#10;
address_ina = 10;
address_inb = 11;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 12;
address_inb = 13;
data_ina = 16'h2;
data_inb = 16'hfffe;
#10;
address_ina = 14;
address_inb = 15;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 16;
address_inb = 17;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 18;
address_inb = 19;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 20;
address_inb = 21;
data_ina = 16'h2;
data_inb = 16'h0;
#10;
address_ina = 22;
address_inb = 23;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 24;
address_inb = 25;
data_ina = 16'hfffe;
data_inb = 16'h0;
#10;
address_ina = 26;
address_inb = 27;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 28;
address_inb = 29;
data_ina = 16'h2;
data_inb = 16'h0;
#10;
address_ina = 30;
address_inb = 31;
data_ina = 16'h0;
data_inb = 16'hfffe;
#10;
address_ina = 32;
address_inb = 33;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 34;
address_inb = 35;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 36;
address_inb = 37;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 38;
address_inb = 39;
data_ina = 16'h2;
data_inb = 16'h0;
#10;
address_ina = 40;
address_inb = 41;
data_ina = 16'hfffe;
data_inb = 16'h0;
#10;
address_ina = 42;
address_inb = 43;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 44;
address_inb = 45;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 46;
address_inb = 47;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 48;
address_inb = 49;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 50;
address_inb = 51;
data_ina = 16'hffff;
data_inb = 16'hfffd;
#10;
address_ina = 52;
address_inb = 53;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 54;
address_inb = 55;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 56;
address_inb = 57;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 58;
address_inb = 59;
data_ina = 16'h0;
data_inb = 16'h2;
#10;
address_ina = 60;
address_inb = 61;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 62;
address_inb = 63;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 64;
address_inb = 65;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 66;
address_inb = 67;
data_ina = 16'hfffe;
data_inb = 16'h0;
#10;
address_ina = 68;
address_inb = 69;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 70;
address_inb = 71;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 72;
address_inb = 73;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 74;
address_inb = 75;
data_ina = 16'h1;
data_inb = 16'h2;
#10;
address_ina = 76;
address_inb = 77;
data_ina = 16'hfffe;
data_inb = 16'h3;
#10;
address_ina = 78;
address_inb = 79;
data_ina = 16'hffff;
data_inb = 16'h2;
#10;
address_ina = 80;
address_inb = 81;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 82;
address_inb = 83;
data_ina = 16'h3;
data_inb = 16'h0;
#10;
address_ina = 84;
address_inb = 85;
data_ina = 16'hffff;
data_inb = 16'hfffe;
#10;
address_ina = 86;
address_inb = 87;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 88;
address_inb = 89;
data_ina = 16'hfffe;
data_inb = 16'hffff;
#10;
address_ina = 90;
address_inb = 91;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 92;
address_inb = 93;
data_ina = 16'hfffe;
data_inb = 16'hfffe;
#10;
address_ina = 94;
address_inb = 95;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 96;
address_inb = 97;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 98;
address_inb = 99;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 100;
address_inb = 101;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 102;
address_inb = 103;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 104;
address_inb = 105;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 106;
address_inb = 107;
data_ina = 16'h0;
data_inb = 16'hfffe;
#10;
address_ina = 108;
address_inb = 109;
data_ina = 16'h1;
data_inb = 16'hfffe;
#10;
address_ina = 110;
address_inb = 111;
data_ina = 16'h2;
data_inb = 16'h2;
#10;
address_ina = 112;
address_inb = 113;
data_ina = 16'hfffe;
data_inb = 16'h0;
#10;
address_ina = 114;
address_inb = 115;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 116;
address_inb = 117;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 118;
address_inb = 119;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 120;
address_inb = 121;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 122;
address_inb = 123;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 124;
address_inb = 125;
data_ina = 16'h0;
data_inb = 16'hfffd;
#10;
address_ina = 126;
address_inb = 127;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 128;
address_inb = 129;
data_ina = 16'h0;
data_inb = 16'hfffe;
#10;
address_ina = 130;
address_inb = 131;
data_ina = 16'hfffd;
data_inb = 16'h0;
#10;
address_ina = 132;
address_inb = 133;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 134;
address_inb = 135;
data_ina = 16'h3;
data_inb = 16'hffff;
#10;
address_ina = 136;
address_inb = 137;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 138;
address_inb = 139;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 140;
address_inb = 141;
data_ina = 16'h1;
data_inb = 16'h2;
#10;
address_ina = 142;
address_inb = 143;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 144;
address_inb = 145;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 146;
address_inb = 147;
data_ina = 16'h2;
data_inb = 16'h1;
#10;
address_ina = 148;
address_inb = 149;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 150;
address_inb = 151;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 152;
address_inb = 153;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 154;
address_inb = 155;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 156;
address_inb = 157;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 158;
address_inb = 159;
data_ina = 16'h1;
data_inb = 16'hfffe;
#10;
address_ina = 160;
address_inb = 161;
data_ina = 16'h1;
data_inb = 16'h2;
#10;
address_ina = 162;
address_inb = 163;
data_ina = 16'hfffe;
data_inb = 16'hffff;
#10;
address_ina = 164;
address_inb = 165;
data_ina = 16'h0;
data_inb = 16'hfffe;
#10;
address_ina = 166;
address_inb = 167;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 168;
address_inb = 169;
data_ina = 16'hfffe;
data_inb = 16'h2;
#10;
address_ina = 170;
address_inb = 171;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 172;
address_inb = 173;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 174;
address_inb = 175;
data_ina = 16'hfffe;
data_inb = 16'h0;
#10;
address_ina = 176;
address_inb = 177;
data_ina = 16'h1;
data_inb = 16'hfffe;
#10;
address_ina = 178;
address_inb = 179;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 180;
address_inb = 181;
data_ina = 16'hfffe;
data_inb = 16'h1;
#10;
address_ina = 182;
address_inb = 183;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 184;
address_inb = 185;
data_ina = 16'h2;
data_inb = 16'h1;
#10;
address_ina = 186;
address_inb = 187;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 188;
address_inb = 189;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 190;
address_inb = 191;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 192;
address_inb = 193;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 194;
address_inb = 195;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 196;
address_inb = 197;
data_ina = 16'h1;
data_inb = 16'hfffe;
#10;
address_ina = 198;
address_inb = 199;
data_ina = 16'hffff;
data_inb = 16'hfffe;
#10;
address_ina = 200;
address_inb = 201;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 202;
address_inb = 203;
data_ina = 16'hffff;
data_inb = 16'h2;
#10;
address_ina = 204;
address_inb = 205;
data_ina = 16'hfffe;
data_inb = 16'h1;
#10;
address_ina = 206;
address_inb = 207;
data_ina = 16'h1;
data_inb = 16'h2;
#10;
address_ina = 208;
address_inb = 209;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 210;
address_inb = 211;
data_ina = 16'h1;
data_inb = 16'hfffe;
#10;
address_ina = 212;
address_inb = 213;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 214;
address_inb = 215;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 216;
address_inb = 217;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 218;
address_inb = 219;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 220;
address_inb = 221;
data_ina = 16'h1;
data_inb = 16'hfffe;
#10;
address_ina = 222;
address_inb = 223;
data_ina = 16'h0;
data_inb = 16'h2;
#10;
address_ina = 224;
address_inb = 225;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 226;
address_inb = 227;
data_ina = 16'hfffe;
data_inb = 16'h1;
#10;
address_ina = 228;
address_inb = 229;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 230;
address_inb = 231;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 232;
address_inb = 233;
data_ina = 16'h0;
data_inb = 16'hfffd;
#10;
address_ina = 234;
address_inb = 235;
data_ina = 16'hffff;
data_inb = 16'hfffd;
#10;
address_ina = 236;
address_inb = 237;
data_ina = 16'hfffe;
data_inb = 16'h1;
#10;
address_ina = 238;
address_inb = 239;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 240;
address_inb = 241;
data_ina = 16'hffff;
data_inb = 16'h2;
#10;
address_ina = 242;
address_inb = 243;
data_ina = 16'hfffe;
data_inb = 16'h1;
#10;
address_ina = 244;
address_inb = 245;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 246;
address_inb = 247;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 248;
address_inb = 249;
data_ina = 16'h2;
data_inb = 16'h1;
#10;
address_ina = 250;
address_inb = 251;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 252;
address_inb = 253;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 254;
address_inb = 255;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
        wait(init_done);
        #30
        we = 0;
        // Start processing
         
		  #38000

        start = 0;



//        wait (wr_req);
//		  wait (!wr_req);
//		   rd_req = 1;
		  wait(done);
		  #20000
rd_req = 1;
        #70 
		  start = 1;
		 #80 
wait(rd_empty)
rd_req = 0;

$display("Finished the NTT test Number %d",test_num);
////Begin test number #70//////////////
rst = 1;

//#1000
start = 1;
mode = 0; //NTT 0 // INTT 1

// Reset for a few clock cycles

#1000

rst = 0;
test_num = test_num + 1;
#1000
we = 1;
address_ina = 0;
address_inb = 1;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 2;
address_inb = 3;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 4;
address_inb = 5;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 6;
address_inb = 7;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 8;
address_inb = 9;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 10;
address_inb = 11;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 12;
address_inb = 13;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 14;
address_inb = 15;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 16;
address_inb = 17;
data_ina = 16'hfffe;
data_inb = 16'h1;
#10;
address_ina = 18;
address_inb = 19;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 20;
address_inb = 21;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 22;
address_inb = 23;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 24;
address_inb = 25;
data_ina = 16'h1;
data_inb = 16'hfffd;
#10;
address_ina = 26;
address_inb = 27;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 28;
address_inb = 29;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 30;
address_inb = 31;
data_ina = 16'hfffe;
data_inb = 16'h3;
#10;
address_ina = 32;
address_inb = 33;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 34;
address_inb = 35;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 36;
address_inb = 37;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 38;
address_inb = 39;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 40;
address_inb = 41;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 42;
address_inb = 43;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 44;
address_inb = 45;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 46;
address_inb = 47;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 48;
address_inb = 49;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 50;
address_inb = 51;
data_ina = 16'h2;
data_inb = 16'hfffe;
#10;
address_ina = 52;
address_inb = 53;
data_ina = 16'hffff;
data_inb = 16'h3;
#10;
address_ina = 54;
address_inb = 55;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 56;
address_inb = 57;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 58;
address_inb = 59;
data_ina = 16'hfffe;
data_inb = 16'h0;
#10;
address_ina = 60;
address_inb = 61;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 62;
address_inb = 63;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 64;
address_inb = 65;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 66;
address_inb = 67;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 68;
address_inb = 69;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 70;
address_inb = 71;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 72;
address_inb = 73;
data_ina = 16'h2;
data_inb = 16'h1;
#10;
address_ina = 74;
address_inb = 75;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 76;
address_inb = 77;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 78;
address_inb = 79;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 80;
address_inb = 81;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 82;
address_inb = 83;
data_ina = 16'h0;
data_inb = 16'hfffd;
#10;
address_ina = 84;
address_inb = 85;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 86;
address_inb = 87;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 88;
address_inb = 89;
data_ina = 16'h2;
data_inb = 16'hffff;
#10;
address_ina = 90;
address_inb = 91;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 92;
address_inb = 93;
data_ina = 16'hfffe;
data_inb = 16'h1;
#10;
address_ina = 94;
address_inb = 95;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 96;
address_inb = 97;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 98;
address_inb = 99;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 100;
address_inb = 101;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 102;
address_inb = 103;
data_ina = 16'hfffe;
data_inb = 16'h2;
#10;
address_ina = 104;
address_inb = 105;
data_ina = 16'h2;
data_inb = 16'h0;
#10;
address_ina = 106;
address_inb = 107;
data_ina = 16'h2;
data_inb = 16'h0;
#10;
address_ina = 108;
address_inb = 109;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 110;
address_inb = 111;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 112;
address_inb = 113;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 114;
address_inb = 115;
data_ina = 16'h0;
data_inb = 16'h3;
#10;
address_ina = 116;
address_inb = 117;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 118;
address_inb = 119;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 120;
address_inb = 121;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 122;
address_inb = 123;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 124;
address_inb = 125;
data_ina = 16'h2;
data_inb = 16'h2;
#10;
address_ina = 126;
address_inb = 127;
data_ina = 16'h0;
data_inb = 16'hfffe;
#10;
address_ina = 128;
address_inb = 129;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 130;
address_inb = 131;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 132;
address_inb = 133;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 134;
address_inb = 135;
data_ina = 16'hfffe;
data_inb = 16'hffff;
#10;
address_ina = 136;
address_inb = 137;
data_ina = 16'h2;
data_inb = 16'h2;
#10;
address_ina = 138;
address_inb = 139;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 140;
address_inb = 141;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 142;
address_inb = 143;
data_ina = 16'h0;
data_inb = 16'h2;
#10;
address_ina = 144;
address_inb = 145;
data_ina = 16'h2;
data_inb = 16'h2;
#10;
address_ina = 146;
address_inb = 147;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 148;
address_inb = 149;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 150;
address_inb = 151;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 152;
address_inb = 153;
data_ina = 16'hfffe;
data_inb = 16'h1;
#10;
address_ina = 154;
address_inb = 155;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 156;
address_inb = 157;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 158;
address_inb = 159;
data_ina = 16'hffff;
data_inb = 16'h2;
#10;
address_ina = 160;
address_inb = 161;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 162;
address_inb = 163;
data_ina = 16'h0;
data_inb = 16'hfffe;
#10;
address_ina = 164;
address_inb = 165;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 166;
address_inb = 167;
data_ina = 16'hfffe;
data_inb = 16'hffff;
#10;
address_ina = 168;
address_inb = 169;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 170;
address_inb = 171;
data_ina = 16'h1;
data_inb = 16'h2;
#10;
address_ina = 172;
address_inb = 173;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 174;
address_inb = 175;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 176;
address_inb = 177;
data_ina = 16'hfffe;
data_inb = 16'h1;
#10;
address_ina = 178;
address_inb = 179;
data_ina = 16'hffff;
data_inb = 16'hfffe;
#10;
address_ina = 180;
address_inb = 181;
data_ina = 16'h2;
data_inb = 16'h0;
#10;
address_ina = 182;
address_inb = 183;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 184;
address_inb = 185;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 186;
address_inb = 187;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 188;
address_inb = 189;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 190;
address_inb = 191;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 192;
address_inb = 193;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 194;
address_inb = 195;
data_ina = 16'h0;
data_inb = 16'hfffe;
#10;
address_ina = 196;
address_inb = 197;
data_ina = 16'h2;
data_inb = 16'h2;
#10;
address_ina = 198;
address_inb = 199;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 200;
address_inb = 201;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 202;
address_inb = 203;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 204;
address_inb = 205;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 206;
address_inb = 207;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 208;
address_inb = 209;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 210;
address_inb = 211;
data_ina = 16'h3;
data_inb = 16'hffff;
#10;
address_ina = 212;
address_inb = 213;
data_ina = 16'h0;
data_inb = 16'hfffe;
#10;
address_ina = 214;
address_inb = 215;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 216;
address_inb = 217;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 218;
address_inb = 219;
data_ina = 16'h3;
data_inb = 16'hffff;
#10;
address_ina = 220;
address_inb = 221;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 222;
address_inb = 223;
data_ina = 16'h2;
data_inb = 16'h2;
#10;
address_ina = 224;
address_inb = 225;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 226;
address_inb = 227;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 228;
address_inb = 229;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 230;
address_inb = 231;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 232;
address_inb = 233;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 234;
address_inb = 235;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 236;
address_inb = 237;
data_ina = 16'h1;
data_inb = 16'h3;
#10;
address_ina = 238;
address_inb = 239;
data_ina = 16'h2;
data_inb = 16'hfffe;
#10;
address_ina = 240;
address_inb = 241;
data_ina = 16'hfffe;
data_inb = 16'h0;
#10;
address_ina = 242;
address_inb = 243;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 244;
address_inb = 245;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 246;
address_inb = 247;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 248;
address_inb = 249;
data_ina = 16'h2;
data_inb = 16'h0;
#10;
address_ina = 250;
address_inb = 251;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 252;
address_inb = 253;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 254;
address_inb = 255;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
        wait(init_done);
        #30
        we = 0;
        // Start processing
         
		  #38000

        start = 0;



//        wait (wr_req);
//		  wait (!wr_req);
//		   rd_req = 1;
		  wait(done);
		  #20000
rd_req = 1;
        #70 
		  start = 1;
		 #80 
wait(rd_empty)
rd_req = 0;

$display("Finished the NTT test Number %d",test_num);
////Begin test number #71//////////////
rst = 1;

//#1000
start = 1;
mode = 0; //NTT 0 // INTT 1

// Reset for a few clock cycles

#1000

rst = 0;
test_num = test_num + 1;
#1000
we = 1;
address_ina = 0;
address_inb = 1;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 2;
address_inb = 3;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 4;
address_inb = 5;
data_ina = 16'h1;
data_inb = 16'hfffe;
#10;
address_ina = 6;
address_inb = 7;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 8;
address_inb = 9;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 10;
address_inb = 11;
data_ina = 16'h2;
data_inb = 16'h0;
#10;
address_ina = 12;
address_inb = 13;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 14;
address_inb = 15;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 16;
address_inb = 17;
data_ina = 16'h2;
data_inb = 16'hffff;
#10;
address_ina = 18;
address_inb = 19;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 20;
address_inb = 21;
data_ina = 16'hfffe;
data_inb = 16'hffff;
#10;
address_ina = 22;
address_inb = 23;
data_ina = 16'h1;
data_inb = 16'h2;
#10;
address_ina = 24;
address_inb = 25;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 26;
address_inb = 27;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 28;
address_inb = 29;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 30;
address_inb = 31;
data_ina = 16'hfffe;
data_inb = 16'h0;
#10;
address_ina = 32;
address_inb = 33;
data_ina = 16'h1;
data_inb = 16'h3;
#10;
address_ina = 34;
address_inb = 35;
data_ina = 16'h1;
data_inb = 16'hfffe;
#10;
address_ina = 36;
address_inb = 37;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 38;
address_inb = 39;
data_ina = 16'hfffe;
data_inb = 16'h2;
#10;
address_ina = 40;
address_inb = 41;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 42;
address_inb = 43;
data_ina = 16'h0;
data_inb = 16'h2;
#10;
address_ina = 44;
address_inb = 45;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 46;
address_inb = 47;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 48;
address_inb = 49;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 50;
address_inb = 51;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 52;
address_inb = 53;
data_ina = 16'hfffe;
data_inb = 16'h1;
#10;
address_ina = 54;
address_inb = 55;
data_ina = 16'h2;
data_inb = 16'hffff;
#10;
address_ina = 56;
address_inb = 57;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 58;
address_inb = 59;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 60;
address_inb = 61;
data_ina = 16'h1;
data_inb = 16'hfffe;
#10;
address_ina = 62;
address_inb = 63;
data_ina = 16'h0;
data_inb = 16'hfffe;
#10;
address_ina = 64;
address_inb = 65;
data_ina = 16'h1;
data_inb = 16'h2;
#10;
address_ina = 66;
address_inb = 67;
data_ina = 16'h2;
data_inb = 16'hffff;
#10;
address_ina = 68;
address_inb = 69;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 70;
address_inb = 71;
data_ina = 16'hffff;
data_inb = 16'hfffe;
#10;
address_ina = 72;
address_inb = 73;
data_ina = 16'h2;
data_inb = 16'h0;
#10;
address_ina = 74;
address_inb = 75;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 76;
address_inb = 77;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 78;
address_inb = 79;
data_ina = 16'hfffe;
data_inb = 16'h0;
#10;
address_ina = 80;
address_inb = 81;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 82;
address_inb = 83;
data_ina = 16'hfffe;
data_inb = 16'h0;
#10;
address_ina = 84;
address_inb = 85;
data_ina = 16'h0;
data_inb = 16'h3;
#10;
address_ina = 86;
address_inb = 87;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 88;
address_inb = 89;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 90;
address_inb = 91;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 92;
address_inb = 93;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 94;
address_inb = 95;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 96;
address_inb = 97;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 98;
address_inb = 99;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 100;
address_inb = 101;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 102;
address_inb = 103;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 104;
address_inb = 105;
data_ina = 16'hffff;
data_inb = 16'hfffe;
#10;
address_ina = 106;
address_inb = 107;
data_ina = 16'h2;
data_inb = 16'h0;
#10;
address_ina = 108;
address_inb = 109;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 110;
address_inb = 111;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 112;
address_inb = 113;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 114;
address_inb = 115;
data_ina = 16'h2;
data_inb = 16'h1;
#10;
address_ina = 116;
address_inb = 117;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 118;
address_inb = 119;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 120;
address_inb = 121;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 122;
address_inb = 123;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 124;
address_inb = 125;
data_ina = 16'hfffe;
data_inb = 16'h0;
#10;
address_ina = 126;
address_inb = 127;
data_ina = 16'h0;
data_inb = 16'hfffd;
#10;
address_ina = 128;
address_inb = 129;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 130;
address_inb = 131;
data_ina = 16'h2;
data_inb = 16'h1;
#10;
address_ina = 132;
address_inb = 133;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 134;
address_inb = 135;
data_ina = 16'hfffe;
data_inb = 16'h0;
#10;
address_ina = 136;
address_inb = 137;
data_ina = 16'h1;
data_inb = 16'h2;
#10;
address_ina = 138;
address_inb = 139;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 140;
address_inb = 141;
data_ina = 16'hfffe;
data_inb = 16'h1;
#10;
address_ina = 142;
address_inb = 143;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 144;
address_inb = 145;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 146;
address_inb = 147;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 148;
address_inb = 149;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 150;
address_inb = 151;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 152;
address_inb = 153;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 154;
address_inb = 155;
data_ina = 16'h1;
data_inb = 16'h2;
#10;
address_ina = 156;
address_inb = 157;
data_ina = 16'h2;
data_inb = 16'h1;
#10;
address_ina = 158;
address_inb = 159;
data_ina = 16'h2;
data_inb = 16'h0;
#10;
address_ina = 160;
address_inb = 161;
data_ina = 16'hffff;
data_inb = 16'h2;
#10;
address_ina = 162;
address_inb = 163;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 164;
address_inb = 165;
data_ina = 16'h1;
data_inb = 16'hfffe;
#10;
address_ina = 166;
address_inb = 167;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 168;
address_inb = 169;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 170;
address_inb = 171;
data_ina = 16'h0;
data_inb = 16'hfffe;
#10;
address_ina = 172;
address_inb = 173;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 174;
address_inb = 175;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 176;
address_inb = 177;
data_ina = 16'hfffe;
data_inb = 16'h1;
#10;
address_ina = 178;
address_inb = 179;
data_ina = 16'h1;
data_inb = 16'h2;
#10;
address_ina = 180;
address_inb = 181;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 182;
address_inb = 183;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 184;
address_inb = 185;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 186;
address_inb = 187;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 188;
address_inb = 189;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 190;
address_inb = 191;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 192;
address_inb = 193;
data_ina = 16'h1;
data_inb = 16'h3;
#10;
address_ina = 194;
address_inb = 195;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 196;
address_inb = 197;
data_ina = 16'hfffd;
data_inb = 16'h2;
#10;
address_ina = 198;
address_inb = 199;
data_ina = 16'h2;
data_inb = 16'h2;
#10;
address_ina = 200;
address_inb = 201;
data_ina = 16'h2;
data_inb = 16'h0;
#10;
address_ina = 202;
address_inb = 203;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 204;
address_inb = 205;
data_ina = 16'h2;
data_inb = 16'hffff;
#10;
address_ina = 206;
address_inb = 207;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 208;
address_inb = 209;
data_ina = 16'hffff;
data_inb = 16'hfffe;
#10;
address_ina = 210;
address_inb = 211;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 212;
address_inb = 213;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 214;
address_inb = 215;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 216;
address_inb = 217;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 218;
address_inb = 219;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 220;
address_inb = 221;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 222;
address_inb = 223;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 224;
address_inb = 225;
data_ina = 16'hfffe;
data_inb = 16'h0;
#10;
address_ina = 226;
address_inb = 227;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 228;
address_inb = 229;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 230;
address_inb = 231;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 232;
address_inb = 233;
data_ina = 16'h2;
data_inb = 16'h0;
#10;
address_ina = 234;
address_inb = 235;
data_ina = 16'h2;
data_inb = 16'hffff;
#10;
address_ina = 236;
address_inb = 237;
data_ina = 16'h2;
data_inb = 16'hffff;
#10;
address_ina = 238;
address_inb = 239;
data_ina = 16'h1;
data_inb = 16'hfffe;
#10;
address_ina = 240;
address_inb = 241;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 242;
address_inb = 243;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 244;
address_inb = 245;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 246;
address_inb = 247;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 248;
address_inb = 249;
data_ina = 16'h1;
data_inb = 16'hfffe;
#10;
address_ina = 250;
address_inb = 251;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 252;
address_inb = 253;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 254;
address_inb = 255;
data_ina = 16'hffff;
data_inb = 16'h3;
#10;
        wait(init_done);
        #30
        we = 0;
        // Start processing
         
		  #38000

        start = 0;



//        wait (wr_req);
//		  wait (!wr_req);
//		   rd_req = 1;
		  wait(done);
		  #20000
rd_req = 1;
        #70 
		  start = 1;
		 #80 
wait(rd_empty)
rd_req = 0;

$display("Finished the NTT test Number %d",test_num);
////Begin test number #72//////////////
rst = 1;

//#1000
start = 1;
mode = 0; //NTT 0 // INTT 1

// Reset for a few clock cycles

#1000

rst = 0;
test_num = test_num + 1;
#1000
we = 1;
address_ina = 0;
address_inb = 1;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 2;
address_inb = 3;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 4;
address_inb = 5;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 6;
address_inb = 7;
data_ina = 16'h2;
data_inb = 16'hffff;
#10;
address_ina = 8;
address_inb = 9;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 10;
address_inb = 11;
data_ina = 16'h1;
data_inb = 16'h2;
#10;
address_ina = 12;
address_inb = 13;
data_ina = 16'h0;
data_inb = 16'hfffd;
#10;
address_ina = 14;
address_inb = 15;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 16;
address_inb = 17;
data_ina = 16'h2;
data_inb = 16'h0;
#10;
address_ina = 18;
address_inb = 19;
data_ina = 16'hfffe;
data_inb = 16'hfffe;
#10;
address_ina = 20;
address_inb = 21;
data_ina = 16'hfffe;
data_inb = 16'h2;
#10;
address_ina = 22;
address_inb = 23;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 24;
address_inb = 25;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 26;
address_inb = 27;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 28;
address_inb = 29;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 30;
address_inb = 31;
data_ina = 16'hffff;
data_inb = 16'hfffe;
#10;
address_ina = 32;
address_inb = 33;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 34;
address_inb = 35;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 36;
address_inb = 37;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 38;
address_inb = 39;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 40;
address_inb = 41;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 42;
address_inb = 43;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 44;
address_inb = 45;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 46;
address_inb = 47;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 48;
address_inb = 49;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 50;
address_inb = 51;
data_ina = 16'h1;
data_inb = 16'hfffe;
#10;
address_ina = 52;
address_inb = 53;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 54;
address_inb = 55;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 56;
address_inb = 57;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 58;
address_inb = 59;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 60;
address_inb = 61;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 62;
address_inb = 63;
data_ina = 16'h2;
data_inb = 16'h0;
#10;
address_ina = 64;
address_inb = 65;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 66;
address_inb = 67;
data_ina = 16'hfffe;
data_inb = 16'h0;
#10;
address_ina = 68;
address_inb = 69;
data_ina = 16'hfffe;
data_inb = 16'h1;
#10;
address_ina = 70;
address_inb = 71;
data_ina = 16'h0;
data_inb = 16'h2;
#10;
address_ina = 72;
address_inb = 73;
data_ina = 16'h2;
data_inb = 16'h1;
#10;
address_ina = 74;
address_inb = 75;
data_ina = 16'h1;
data_inb = 16'h2;
#10;
address_ina = 76;
address_inb = 77;
data_ina = 16'hfffe;
data_inb = 16'hffff;
#10;
address_ina = 78;
address_inb = 79;
data_ina = 16'h1;
data_inb = 16'hfffe;
#10;
address_ina = 80;
address_inb = 81;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 82;
address_inb = 83;
data_ina = 16'hfffd;
data_inb = 16'h1;
#10;
address_ina = 84;
address_inb = 85;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 86;
address_inb = 87;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 88;
address_inb = 89;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 90;
address_inb = 91;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 92;
address_inb = 93;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 94;
address_inb = 95;
data_ina = 16'h0;
data_inb = 16'hfffe;
#10;
address_ina = 96;
address_inb = 97;
data_ina = 16'hfffe;
data_inb = 16'h2;
#10;
address_ina = 98;
address_inb = 99;
data_ina = 16'h0;
data_inb = 16'h2;
#10;
address_ina = 100;
address_inb = 101;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 102;
address_inb = 103;
data_ina = 16'h0;
data_inb = 16'hfffe;
#10;
address_ina = 104;
address_inb = 105;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 106;
address_inb = 107;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 108;
address_inb = 109;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 110;
address_inb = 111;
data_ina = 16'hfffe;
data_inb = 16'hfffe;
#10;
address_ina = 112;
address_inb = 113;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 114;
address_inb = 115;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 116;
address_inb = 117;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 118;
address_inb = 119;
data_ina = 16'hffff;
data_inb = 16'h2;
#10;
address_ina = 120;
address_inb = 121;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 122;
address_inb = 123;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 124;
address_inb = 125;
data_ina = 16'h2;
data_inb = 16'h0;
#10;
address_ina = 126;
address_inb = 127;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 128;
address_inb = 129;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 130;
address_inb = 131;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 132;
address_inb = 133;
data_ina = 16'h0;
data_inb = 16'h2;
#10;
address_ina = 134;
address_inb = 135;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 136;
address_inb = 137;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 138;
address_inb = 139;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 140;
address_inb = 141;
data_ina = 16'hfffe;
data_inb = 16'hffff;
#10;
address_ina = 142;
address_inb = 143;
data_ina = 16'hfffe;
data_inb = 16'h0;
#10;
address_ina = 144;
address_inb = 145;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 146;
address_inb = 147;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 148;
address_inb = 149;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 150;
address_inb = 151;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 152;
address_inb = 153;
data_ina = 16'h2;
data_inb = 16'hffff;
#10;
address_ina = 154;
address_inb = 155;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 156;
address_inb = 157;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 158;
address_inb = 159;
data_ina = 16'hffff;
data_inb = 16'h2;
#10;
address_ina = 160;
address_inb = 161;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 162;
address_inb = 163;
data_ina = 16'hfffe;
data_inb = 16'h0;
#10;
address_ina = 164;
address_inb = 165;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 166;
address_inb = 167;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 168;
address_inb = 169;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 170;
address_inb = 171;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 172;
address_inb = 173;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 174;
address_inb = 175;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 176;
address_inb = 177;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 178;
address_inb = 179;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 180;
address_inb = 181;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 182;
address_inb = 183;
data_ina = 16'h0;
data_inb = 16'h2;
#10;
address_ina = 184;
address_inb = 185;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 186;
address_inb = 187;
data_ina = 16'h0;
data_inb = 16'hfffe;
#10;
address_ina = 188;
address_inb = 189;
data_ina = 16'h1;
data_inb = 16'hfffe;
#10;
address_ina = 190;
address_inb = 191;
data_ina = 16'h2;
data_inb = 16'hffff;
#10;
address_ina = 192;
address_inb = 193;
data_ina = 16'hffff;
data_inb = 16'h2;
#10;
address_ina = 194;
address_inb = 195;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 196;
address_inb = 197;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 198;
address_inb = 199;
data_ina = 16'h2;
data_inb = 16'h1;
#10;
address_ina = 200;
address_inb = 201;
data_ina = 16'hfffe;
data_inb = 16'h0;
#10;
address_ina = 202;
address_inb = 203;
data_ina = 16'h2;
data_inb = 16'hffff;
#10;
address_ina = 204;
address_inb = 205;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 206;
address_inb = 207;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 208;
address_inb = 209;
data_ina = 16'h0;
data_inb = 16'h2;
#10;
address_ina = 210;
address_inb = 211;
data_ina = 16'h2;
data_inb = 16'h0;
#10;
address_ina = 212;
address_inb = 213;
data_ina = 16'h1;
data_inb = 16'hfffe;
#10;
address_ina = 214;
address_inb = 215;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 216;
address_inb = 217;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 218;
address_inb = 219;
data_ina = 16'h0;
data_inb = 16'h2;
#10;
address_ina = 220;
address_inb = 221;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 222;
address_inb = 223;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 224;
address_inb = 225;
data_ina = 16'h2;
data_inb = 16'hfffe;
#10;
address_ina = 226;
address_inb = 227;
data_ina = 16'h2;
data_inb = 16'h0;
#10;
address_ina = 228;
address_inb = 229;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 230;
address_inb = 231;
data_ina = 16'h1;
data_inb = 16'h2;
#10;
address_ina = 232;
address_inb = 233;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 234;
address_inb = 235;
data_ina = 16'h3;
data_inb = 16'hffff;
#10;
address_ina = 236;
address_inb = 237;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 238;
address_inb = 239;
data_ina = 16'hffff;
data_inb = 16'hfffe;
#10;
address_ina = 240;
address_inb = 241;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 242;
address_inb = 243;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 244;
address_inb = 245;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 246;
address_inb = 247;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 248;
address_inb = 249;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 250;
address_inb = 251;
data_ina = 16'hfffe;
data_inb = 16'h0;
#10;
address_ina = 252;
address_inb = 253;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 254;
address_inb = 255;
data_ina = 16'h0;
data_inb = 16'hfffe;
#10;
        wait(init_done);
        #30
        we = 0;
        // Start processing
         
		  #38000

        start = 0;



//        wait (wr_req);
//		  wait (!wr_req);
//		   rd_req = 1;
		  wait(done);
		  #20000
rd_req = 1;
        #70 
		  start = 1;
		 #80 
wait(rd_empty)
rd_req = 0;

$display("Finished the NTT test Number %d",test_num);
////Begin test number #73//////////////
rst = 1;

//#1000
start = 1;
mode = 0; //NTT 0 // INTT 1

// Reset for a few clock cycles

#1000

rst = 0;
test_num = test_num + 1;
#1000
we = 1;
address_ina = 0;
address_inb = 1;
data_ina = 16'hffff;
data_inb = 16'hfffe;
#10;
address_ina = 2;
address_inb = 3;
data_ina = 16'h1;
data_inb = 16'h2;
#10;
address_ina = 4;
address_inb = 5;
data_ina = 16'h0;
data_inb = 16'h2;
#10;
address_ina = 6;
address_inb = 7;
data_ina = 16'hfffe;
data_inb = 16'hfffe;
#10;
address_ina = 8;
address_inb = 9;
data_ina = 16'h1;
data_inb = 16'h2;
#10;
address_ina = 10;
address_inb = 11;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 12;
address_inb = 13;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 14;
address_inb = 15;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 16;
address_inb = 17;
data_ina = 16'h3;
data_inb = 16'h0;
#10;
address_ina = 18;
address_inb = 19;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 20;
address_inb = 21;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 22;
address_inb = 23;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 24;
address_inb = 25;
data_ina = 16'h2;
data_inb = 16'h1;
#10;
address_ina = 26;
address_inb = 27;
data_ina = 16'hfffe;
data_inb = 16'hffff;
#10;
address_ina = 28;
address_inb = 29;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 30;
address_inb = 31;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 32;
address_inb = 33;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 34;
address_inb = 35;
data_ina = 16'hfffe;
data_inb = 16'hfffe;
#10;
address_ina = 36;
address_inb = 37;
data_ina = 16'h2;
data_inb = 16'h0;
#10;
address_ina = 38;
address_inb = 39;
data_ina = 16'h2;
data_inb = 16'hffff;
#10;
address_ina = 40;
address_inb = 41;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 42;
address_inb = 43;
data_ina = 16'h2;
data_inb = 16'hfffe;
#10;
address_ina = 44;
address_inb = 45;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 46;
address_inb = 47;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 48;
address_inb = 49;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 50;
address_inb = 51;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 52;
address_inb = 53;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 54;
address_inb = 55;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 56;
address_inb = 57;
data_ina = 16'hffff;
data_inb = 16'hfffe;
#10;
address_ina = 58;
address_inb = 59;
data_ina = 16'hffff;
data_inb = 16'h2;
#10;
address_ina = 60;
address_inb = 61;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 62;
address_inb = 63;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 64;
address_inb = 65;
data_ina = 16'h0;
data_inb = 16'hfffe;
#10;
address_ina = 66;
address_inb = 67;
data_ina = 16'hfffd;
data_inb = 16'h1;
#10;
address_ina = 68;
address_inb = 69;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 70;
address_inb = 71;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 72;
address_inb = 73;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 74;
address_inb = 75;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 76;
address_inb = 77;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 78;
address_inb = 79;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 80;
address_inb = 81;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 82;
address_inb = 83;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 84;
address_inb = 85;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 86;
address_inb = 87;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 88;
address_inb = 89;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 90;
address_inb = 91;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 92;
address_inb = 93;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 94;
address_inb = 95;
data_ina = 16'h1;
data_inb = 16'h2;
#10;
address_ina = 96;
address_inb = 97;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 98;
address_inb = 99;
data_ina = 16'h0;
data_inb = 16'h2;
#10;
address_ina = 100;
address_inb = 101;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 102;
address_inb = 103;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 104;
address_inb = 105;
data_ina = 16'hfffe;
data_inb = 16'hfffe;
#10;
address_ina = 106;
address_inb = 107;
data_ina = 16'h2;
data_inb = 16'h1;
#10;
address_ina = 108;
address_inb = 109;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 110;
address_inb = 111;
data_ina = 16'hfffe;
data_inb = 16'hfffd;
#10;
address_ina = 112;
address_inb = 113;
data_ina = 16'h0;
data_inb = 16'h2;
#10;
address_ina = 114;
address_inb = 115;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 116;
address_inb = 117;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 118;
address_inb = 119;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 120;
address_inb = 121;
data_ina = 16'hfffe;
data_inb = 16'h0;
#10;
address_ina = 122;
address_inb = 123;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 124;
address_inb = 125;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 126;
address_inb = 127;
data_ina = 16'h2;
data_inb = 16'hffff;
#10;
address_ina = 128;
address_inb = 129;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 130;
address_inb = 131;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 132;
address_inb = 133;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 134;
address_inb = 135;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 136;
address_inb = 137;
data_ina = 16'hfffd;
data_inb = 16'h1;
#10;
address_ina = 138;
address_inb = 139;
data_ina = 16'hfffe;
data_inb = 16'h1;
#10;
address_ina = 140;
address_inb = 141;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 142;
address_inb = 143;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 144;
address_inb = 145;
data_ina = 16'h1;
data_inb = 16'h2;
#10;
address_ina = 146;
address_inb = 147;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 148;
address_inb = 149;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 150;
address_inb = 151;
data_ina = 16'h2;
data_inb = 16'h0;
#10;
address_ina = 152;
address_inb = 153;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 154;
address_inb = 155;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 156;
address_inb = 157;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 158;
address_inb = 159;
data_ina = 16'h0;
data_inb = 16'hfffe;
#10;
address_ina = 160;
address_inb = 161;
data_ina = 16'hfffe;
data_inb = 16'h0;
#10;
address_ina = 162;
address_inb = 163;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 164;
address_inb = 165;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 166;
address_inb = 167;
data_ina = 16'h0;
data_inb = 16'hfffe;
#10;
address_ina = 168;
address_inb = 169;
data_ina = 16'h0;
data_inb = 16'h2;
#10;
address_ina = 170;
address_inb = 171;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 172;
address_inb = 173;
data_ina = 16'h2;
data_inb = 16'h1;
#10;
address_ina = 174;
address_inb = 175;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 176;
address_inb = 177;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 178;
address_inb = 179;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 180;
address_inb = 181;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 182;
address_inb = 183;
data_ina = 16'h2;
data_inb = 16'hffff;
#10;
address_ina = 184;
address_inb = 185;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 186;
address_inb = 187;
data_ina = 16'h3;
data_inb = 16'h0;
#10;
address_ina = 188;
address_inb = 189;
data_ina = 16'h0;
data_inb = 16'hfffe;
#10;
address_ina = 190;
address_inb = 191;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 192;
address_inb = 193;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 194;
address_inb = 195;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 196;
address_inb = 197;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 198;
address_inb = 199;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 200;
address_inb = 201;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 202;
address_inb = 203;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 204;
address_inb = 205;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 206;
address_inb = 207;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 208;
address_inb = 209;
data_ina = 16'hfffe;
data_inb = 16'h1;
#10;
address_ina = 210;
address_inb = 211;
data_ina = 16'hfffe;
data_inb = 16'hffff;
#10;
address_ina = 212;
address_inb = 213;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 214;
address_inb = 215;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 216;
address_inb = 217;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 218;
address_inb = 219;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 220;
address_inb = 221;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 222;
address_inb = 223;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 224;
address_inb = 225;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 226;
address_inb = 227;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 228;
address_inb = 229;
data_ina = 16'h0;
data_inb = 16'h3;
#10;
address_ina = 230;
address_inb = 231;
data_ina = 16'hfffe;
data_inb = 16'h1;
#10;
address_ina = 232;
address_inb = 233;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 234;
address_inb = 235;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 236;
address_inb = 237;
data_ina = 16'h2;
data_inb = 16'h0;
#10;
address_ina = 238;
address_inb = 239;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 240;
address_inb = 241;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 242;
address_inb = 243;
data_ina = 16'h1;
data_inb = 16'h2;
#10;
address_ina = 244;
address_inb = 245;
data_ina = 16'h2;
data_inb = 16'h1;
#10;
address_ina = 246;
address_inb = 247;
data_ina = 16'h2;
data_inb = 16'h2;
#10;
address_ina = 248;
address_inb = 249;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 250;
address_inb = 251;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 252;
address_inb = 253;
data_ina = 16'h3;
data_inb = 16'h1;
#10;
address_ina = 254;
address_inb = 255;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
        wait(init_done);
        #30
        we = 0;
        // Start processing
         
		  #38000

        start = 0;



//        wait (wr_req);
//		  wait (!wr_req);
//		   rd_req = 1;
		  wait(done);
		  #20000
rd_req = 1;
        #70 
		  start = 1;
		 #80 
wait(rd_empty)
rd_req = 0;

$display("Finished the NTT test Number %d",test_num);
////Begin test number #79//////////////
rst = 1;

//#1000
start = 1;
mode = 1; //NTT 0 // INTT 1

// Reset for a few clock cycles

#1000

rst = 0;
test_num = test_num + 1;
#1000
we = 1;
address_ina = 0;
address_inb = 1;
data_ina = 16'h5b;
data_inb = 16'h275;
#10;
address_ina = 2;
address_inb = 3;
data_ina = 16'hffe6;
data_inb = 16'hfe2d;
#10;
address_ina = 4;
address_inb = 5;
data_ina = 16'hfc29;
data_inb = 16'hfe3f;
#10;
address_ina = 6;
address_inb = 7;
data_ina = 16'hfc8f;
data_inb = 16'h58b;
#10;
address_ina = 8;
address_inb = 9;
data_ina = 16'hfef6;
data_inb = 16'hfd5c;
#10;
address_ina = 10;
address_inb = 11;
data_ina = 16'hfff2;
data_inb = 16'hfb87;
#10;
address_ina = 12;
address_inb = 13;
data_ina = 16'h19a;
data_inb = 16'hfb8c;
#10;
address_ina = 14;
address_inb = 15;
data_ina = 16'h3d6;
data_inb = 16'h4b9;
#10;
address_ina = 16;
address_inb = 17;
data_ina = 16'hfed2;
data_inb = 16'h43b;
#10;
address_ina = 18;
address_inb = 19;
data_ina = 16'hfaf3;
data_inb = 16'hfd7f;
#10;
address_ina = 20;
address_inb = 21;
data_ina = 16'hff12;
data_inb = 16'hfff0;
#10;
address_ina = 22;
address_inb = 23;
data_ina = 16'hfe0d;
data_inb = 16'hfbbc;
#10;
address_ina = 24;
address_inb = 25;
data_ina = 16'h5b6;
data_inb = 16'hfa32;
#10;
address_ina = 26;
address_inb = 27;
data_ina = 16'hfad9;
data_inb = 16'hfb2d;
#10;
address_ina = 28;
address_inb = 29;
data_ina = 16'hffc2;
data_inb = 16'h656;
#10;
address_ina = 30;
address_inb = 31;
data_ina = 16'hff7f;
data_inb = 16'hfcf1;
#10;
address_ina = 32;
address_inb = 33;
data_ina = 16'h1f3;
data_inb = 16'hff12;
#10;
address_ina = 34;
address_inb = 35;
data_ina = 16'hfbde;
data_inb = 16'hfc6f;
#10;
address_ina = 36;
address_inb = 37;
data_ina = 16'h66b;
data_inb = 16'hfbde;
#10;
address_ina = 38;
address_inb = 39;
data_ina = 16'h14b;
data_inb = 16'hff85;
#10;
address_ina = 40;
address_inb = 41;
data_ina = 16'hf9c3;
data_inb = 16'h3ae;
#10;
address_ina = 42;
address_inb = 43;
data_ina = 16'hfdf5;
data_inb = 16'h297;
#10;
address_ina = 44;
address_inb = 45;
data_ina = 16'hfcb7;
data_inb = 16'h65;
#10;
address_ina = 46;
address_inb = 47;
data_ina = 16'h304;
data_inb = 16'h60c;
#10;
address_ina = 48;
address_inb = 49;
data_ina = 16'hff1c;
data_inb = 16'h643;
#10;
address_ina = 50;
address_inb = 51;
data_ina = 16'h1a4;
data_inb = 16'hfd1f;
#10;
address_ina = 52;
address_inb = 53;
data_ina = 16'hfbc4;
data_inb = 16'h5f4;
#10;
address_ina = 54;
address_inb = 55;
data_ina = 16'hfa25;
data_inb = 16'h4ae;
#10;
address_ina = 56;
address_inb = 57;
data_ina = 16'h603;
data_inb = 16'h42b;
#10;
address_ina = 58;
address_inb = 59;
data_ina = 16'h47;
data_inb = 16'h26f;
#10;
address_ina = 60;
address_inb = 61;
data_ina = 16'hfba8;
data_inb = 16'hfdd1;
#10;
address_ina = 62;
address_inb = 63;
data_ina = 16'hfd64;
data_inb = 16'hfe83;
#10;
address_ina = 64;
address_inb = 65;
data_ina = 16'hffbb;
data_inb = 16'h62;
#10;
address_ina = 66;
address_inb = 67;
data_ina = 16'h9;
data_inb = 16'hfa72;
#10;
address_ina = 68;
address_inb = 69;
data_ina = 16'hff0f;
data_inb = 16'hf9bb;
#10;
address_ina = 70;
address_inb = 71;
data_ina = 16'h56c;
data_inb = 16'h594;
#10;
address_ina = 72;
address_inb = 73;
data_ina = 16'h46d;
data_inb = 16'h480;
#10;
address_ina = 74;
address_inb = 75;
data_ina = 16'h11b;
data_inb = 16'hfe40;
#10;
address_ina = 76;
address_inb = 77;
data_ina = 16'ha1;
data_inb = 16'hfff5;
#10;
address_ina = 78;
address_inb = 79;
data_ina = 16'hff0d;
data_inb = 16'hff79;
#10;
address_ina = 80;
address_inb = 81;
data_ina = 16'h40f;
data_inb = 16'h36f;
#10;
address_ina = 82;
address_inb = 83;
data_ina = 16'h28b;
data_inb = 16'h2b7;
#10;
address_ina = 84;
address_inb = 85;
data_ina = 16'h406;
data_inb = 16'h10e;
#10;
address_ina = 86;
address_inb = 87;
data_ina = 16'hffe9;
data_inb = 16'h4e1;
#10;
address_ina = 88;
address_inb = 89;
data_ina = 16'hfcf4;
data_inb = 16'h5f2;
#10;
address_ina = 90;
address_inb = 91;
data_ina = 16'h11;
data_inb = 16'h38d;
#10;
address_ina = 92;
address_inb = 93;
data_ina = 16'hff70;
data_inb = 16'h563;
#10;
address_ina = 94;
address_inb = 95;
data_ina = 16'h4b2;
data_inb = 16'hff57;
#10;
address_ina = 96;
address_inb = 97;
data_ina = 16'hfe68;
data_inb = 16'h3de;
#10;
address_ina = 98;
address_inb = 99;
data_ina = 16'hfb42;
data_inb = 16'hf9be;
#10;
address_ina = 100;
address_inb = 101;
data_ina = 16'hfec3;
data_inb = 16'hfb48;
#10;
address_ina = 102;
address_inb = 103;
data_ina = 16'hfe0f;
data_inb = 16'h226;
#10;
address_ina = 104;
address_inb = 105;
data_ina = 16'h2a9;
data_inb = 16'h472;
#10;
address_ina = 106;
address_inb = 107;
data_ina = 16'hfe02;
data_inb = 16'hf9;
#10;
address_ina = 108;
address_inb = 109;
data_ina = 16'h3d5;
data_inb = 16'hfda2;
#10;
address_ina = 110;
address_inb = 111;
data_ina = 16'h444;
data_inb = 16'hff76;
#10;
address_ina = 112;
address_inb = 113;
data_ina = 16'hb5;
data_inb = 16'h168;
#10;
address_ina = 114;
address_inb = 115;
data_ina = 16'h676;
data_inb = 16'hfa37;
#10;
address_ina = 116;
address_inb = 117;
data_ina = 16'hfddc;
data_inb = 16'hfa29;
#10;
address_ina = 118;
address_inb = 119;
data_ina = 16'hfaae;
data_inb = 16'hfe3d;
#10;
address_ina = 120;
address_inb = 121;
data_ina = 16'h1dd;
data_inb = 16'hfc07;
#10;
address_ina = 122;
address_inb = 123;
data_ina = 16'hffea;
data_inb = 16'hff5b;
#10;
address_ina = 124;
address_inb = 125;
data_ina = 16'h59b;
data_inb = 16'h512;
#10;
address_ina = 126;
address_inb = 127;
data_ina = 16'hfdaa;
data_inb = 16'hfab4;
#10;
address_ina = 128;
address_inb = 129;
data_ina = 16'hf9d1;
data_inb = 16'hfdab;
#10;
address_ina = 130;
address_inb = 131;
data_ina = 16'h3bf;
data_inb = 16'h455;
#10;
address_ina = 132;
address_inb = 133;
data_ina = 16'hfd20;
data_inb = 16'hfdc7;
#10;
address_ina = 134;
address_inb = 135;
data_ina = 16'h553;
data_inb = 16'h3d7;
#10;
address_ina = 136;
address_inb = 137;
data_ina = 16'hfd72;
data_inb = 16'hfc7b;
#10;
address_ina = 138;
address_inb = 139;
data_ina = 16'hfccc;
data_inb = 16'hfff6;
#10;
address_ina = 140;
address_inb = 141;
data_ina = 16'h2b;
data_inb = 16'h8c;
#10;
address_ina = 142;
address_inb = 143;
data_ina = 16'h2d4;
data_inb = 16'h300;
#10;
address_ina = 144;
address_inb = 145;
data_ina = 16'h254;
data_inb = 16'hfe53;
#10;
address_ina = 146;
address_inb = 147;
data_ina = 16'hfa89;
data_inb = 16'hf996;
#10;
address_ina = 148;
address_inb = 149;
data_ina = 16'h540;
data_inb = 16'hfaf0;
#10;
address_ina = 150;
address_inb = 151;
data_ina = 16'hfe8e;
data_inb = 16'h625;
#10;
address_ina = 152;
address_inb = 153;
data_ina = 16'hd1;
data_inb = 16'h48d;
#10;
address_ina = 154;
address_inb = 155;
data_ina = 16'hfe01;
data_inb = 16'h663;
#10;
address_ina = 156;
address_inb = 157;
data_ina = 16'hfe55;
data_inb = 16'hfa28;
#10;
address_ina = 158;
address_inb = 159;
data_ina = 16'h3ee;
data_inb = 16'h201;
#10;
address_ina = 160;
address_inb = 161;
data_ina = 16'hfdb8;
data_inb = 16'hfdc1;
#10;
address_ina = 162;
address_inb = 163;
data_ina = 16'h5f2;
data_inb = 16'h419;
#10;
address_ina = 164;
address_inb = 165;
data_ina = 16'h2ee;
data_inb = 16'h645;
#10;
address_ina = 166;
address_inb = 167;
data_ina = 16'hd2;
data_inb = 16'h367;
#10;
address_ina = 168;
address_inb = 169;
data_ina = 16'h2bb;
data_inb = 16'hfd3e;
#10;
address_ina = 170;
address_inb = 171;
data_ina = 16'hf9d8;
data_inb = 16'hfa5a;
#10;
address_ina = 172;
address_inb = 173;
data_ina = 16'h502;
data_inb = 16'hfbc3;
#10;
address_ina = 174;
address_inb = 175;
data_ina = 16'hfe07;
data_inb = 16'h2c9;
#10;
address_ina = 176;
address_inb = 177;
data_ina = 16'hfbac;
data_inb = 16'h27d;
#10;
address_ina = 178;
address_inb = 179;
data_ina = 16'hfd18;
data_inb = 16'h394;
#10;
address_ina = 180;
address_inb = 181;
data_ina = 16'h123;
data_inb = 16'h26b;
#10;
address_ina = 182;
address_inb = 183;
data_ina = 16'h6e;
data_inb = 16'hfea8;
#10;
address_ina = 184;
address_inb = 185;
data_ina = 16'h159;
data_inb = 16'hfec7;
#10;
address_ina = 186;
address_inb = 187;
data_ina = 16'h517;
data_inb = 16'h3dd;
#10;
address_ina = 188;
address_inb = 189;
data_ina = 16'hfcff;
data_inb = 16'h3d9;
#10;
address_ina = 190;
address_inb = 191;
data_ina = 16'h216;
data_inb = 16'h378;
#10;
address_ina = 192;
address_inb = 193;
data_ina = 16'hfe17;
data_inb = 16'hfa9e;
#10;
address_ina = 194;
address_inb = 195;
data_ina = 16'hfdbf;
data_inb = 16'hfc71;
#10;
address_ina = 196;
address_inb = 197;
data_ina = 16'hfd16;
data_inb = 16'hfeaa;
#10;
address_ina = 198;
address_inb = 199;
data_ina = 16'h98;
data_inb = 16'hfb58;
#10;
address_ina = 200;
address_inb = 201;
data_ina = 16'h36b;
data_inb = 16'hfd52;
#10;
address_ina = 202;
address_inb = 203;
data_ina = 16'h449;
data_inb = 16'h515;
#10;
address_ina = 204;
address_inb = 205;
data_ina = 16'hfcc1;
data_inb = 16'h19b;
#10;
address_ina = 206;
address_inb = 207;
data_ina = 16'hfd87;
data_inb = 16'hc2;
#10;
address_ina = 208;
address_inb = 209;
data_ina = 16'hff04;
data_inb = 16'hfcde;
#10;
address_ina = 210;
address_inb = 211;
data_ina = 16'hfab3;
data_inb = 16'hfcb2;
#10;
address_ina = 212;
address_inb = 213;
data_ina = 16'hfdd9;
data_inb = 16'hfbda;
#10;
address_ina = 214;
address_inb = 215;
data_ina = 16'hfae5;
data_inb = 16'h221;
#10;
address_ina = 216;
address_inb = 217;
data_ina = 16'h308;
data_inb = 16'hfd16;
#10;
address_ina = 218;
address_inb = 219;
data_ina = 16'h23;
data_inb = 16'h1ce;
#10;
address_ina = 220;
address_inb = 221;
data_ina = 16'h1be;
data_inb = 16'h29f;
#10;
address_ina = 222;
address_inb = 223;
data_ina = 16'hfd5c;
data_inb = 16'hfbe8;
#10;
address_ina = 224;
address_inb = 225;
data_ina = 16'h1ec;
data_inb = 16'hf9a9;
#10;
address_ina = 226;
address_inb = 227;
data_ina = 16'hfe65;
data_inb = 16'hfdc5;
#10;
address_ina = 228;
address_inb = 229;
data_ina = 16'h405;
data_inb = 16'hff86;
#10;
address_ina = 230;
address_inb = 231;
data_ina = 16'h4b1;
data_inb = 16'hfa5c;
#10;
address_ina = 232;
address_inb = 233;
data_ina = 16'h5f5;
data_inb = 16'h443;
#10;
address_ina = 234;
address_inb = 235;
data_ina = 16'hfcbe;
data_inb = 16'h12a;
#10;
address_ina = 236;
address_inb = 237;
data_ina = 16'h60c;
data_inb = 16'hfd19;
#10;
address_ina = 238;
address_inb = 239;
data_ina = 16'h8b;
data_inb = 16'hf9df;
#10;
address_ina = 240;
address_inb = 241;
data_ina = 16'hfef7;
data_inb = 16'ha3;
#10;
address_ina = 242;
address_inb = 243;
data_ina = 16'hfad7;
data_inb = 16'h3b4;
#10;
address_ina = 244;
address_inb = 245;
data_ina = 16'hfce3;
data_inb = 16'hfb58;
#10;
address_ina = 246;
address_inb = 247;
data_ina = 16'h509;
data_inb = 16'h46f;
#10;
address_ina = 248;
address_inb = 249;
data_ina = 16'hfa85;
data_inb = 16'hff71;
#10;
address_ina = 250;
address_inb = 251;
data_ina = 16'h25c;
data_inb = 16'h224;
#10;
address_ina = 252;
address_inb = 253;
data_ina = 16'hfe62;
data_inb = 16'h2ed;
#10;
address_ina = 254;
address_inb = 255;
data_ina = 16'hfd66;
data_inb = 16'hffd8;
#10;
        wait(init_done);
        #30
        we = 0;
        // Start processing
         
		  #38000

        start = 0;



//        wait (wr_req);
//		  wait (!wr_req);
//		   rd_req = 1;
		  wait(done);
		  #20000
rd_req = 1;
        #70 
		  start = 1;
		 #80 
wait(rd_empty)
rd_req = 0;

$display("Finished the NTT test Number %d",test_num);
////Begin test number #75//////////////
rst = 1;

//#1000
start = 1;
mode = 1; //NTT 0 // INTT 1

// Reset for a few clock cycles

#1000

rst = 0;
test_num = test_num + 1;
#1000
we = 1;
address_ina = 0;
address_inb = 1;
data_ina = 16'hfb85;
data_inb = 16'hfe5d;
#10;
address_ina = 2;
address_inb = 3;
data_ina = 16'hff39;
data_inb = 16'h5db;
#10;
address_ina = 4;
address_inb = 5;
data_ina = 16'h48;
data_inb = 16'h162;
#10;
address_ina = 6;
address_inb = 7;
data_ina = 16'hfcc1;
data_inb = 16'hfeac;
#10;
address_ina = 8;
address_inb = 9;
data_ina = 16'h80;
data_inb = 16'hfe18;
#10;
address_ina = 10;
address_inb = 11;
data_ina = 16'h4e4;
data_inb = 16'hfa72;
#10;
address_ina = 12;
address_inb = 13;
data_ina = 16'h7f;
data_inb = 16'hfdc1;
#10;
address_ina = 14;
address_inb = 15;
data_ina = 16'h1aa;
data_inb = 16'hfb18;
#10;
address_ina = 16;
address_inb = 17;
data_ina = 16'h54a;
data_inb = 16'h104;
#10;
address_ina = 18;
address_inb = 19;
data_ina = 16'hfad9;
data_inb = 16'h4c8;
#10;
address_ina = 20;
address_inb = 21;
data_ina = 16'hfaca;
data_inb = 16'hffd5;
#10;
address_ina = 22;
address_inb = 23;
data_ina = 16'hfb22;
data_inb = 16'h23c;
#10;
address_ina = 24;
address_inb = 25;
data_ina = 16'h15c;
data_inb = 16'hfb18;
#10;
address_ina = 26;
address_inb = 27;
data_ina = 16'hfe5b;
data_inb = 16'hf9cb;
#10;
address_ina = 28;
address_inb = 29;
data_ina = 16'hfaea;
data_inb = 16'h33;
#10;
address_ina = 30;
address_inb = 31;
data_ina = 16'hfe00;
data_inb = 16'hfe54;
#10;
address_ina = 32;
address_inb = 33;
data_ina = 16'h43f;
data_inb = 16'hfc71;
#10;
address_ina = 34;
address_inb = 35;
data_ina = 16'hffcc;
data_inb = 16'hfd12;
#10;
address_ina = 36;
address_inb = 37;
data_ina = 16'hfee4;
data_inb = 16'h3ef;
#10;
address_ina = 38;
address_inb = 39;
data_ina = 16'h1a3;
data_inb = 16'h224;
#10;
address_ina = 40;
address_inb = 41;
data_ina = 16'h106;
data_inb = 16'hff50;
#10;
address_ina = 42;
address_inb = 43;
data_ina = 16'h554;
data_inb = 16'hfe0e;
#10;
address_ina = 44;
address_inb = 45;
data_ina = 16'hfbf1;
data_inb = 16'h5f8;
#10;
address_ina = 46;
address_inb = 47;
data_ina = 16'h648;
data_inb = 16'h1c1;
#10;
address_ina = 48;
address_inb = 49;
data_ina = 16'h49e;
data_inb = 16'h23c;
#10;
address_ina = 50;
address_inb = 51;
data_ina = 16'h164;
data_inb = 16'hfbda;
#10;
address_ina = 52;
address_inb = 53;
data_ina = 16'hfe71;
data_inb = 16'h54d;
#10;
address_ina = 54;
address_inb = 55;
data_ina = 16'hfd03;
data_inb = 16'h19e;
#10;
address_ina = 56;
address_inb = 57;
data_ina = 16'h5da;
data_inb = 16'hfc84;
#10;
address_ina = 58;
address_inb = 59;
data_ina = 16'hfb57;
data_inb = 16'h4da;
#10;
address_ina = 60;
address_inb = 61;
data_ina = 16'hfe7f;
data_inb = 16'hfd46;
#10;
address_ina = 62;
address_inb = 63;
data_ina = 16'hfe19;
data_inb = 16'hb8;
#10;
address_ina = 64;
address_inb = 65;
data_ina = 16'hfdd7;
data_inb = 16'h277;
#10;
address_ina = 66;
address_inb = 67;
data_ina = 16'h564;
data_inb = 16'hfd59;
#10;
address_ina = 68;
address_inb = 69;
data_ina = 16'hfc88;
data_inb = 16'hfc51;
#10;
address_ina = 70;
address_inb = 71;
data_ina = 16'h1e4;
data_inb = 16'h1d2;
#10;
address_ina = 72;
address_inb = 73;
data_ina = 16'hfce3;
data_inb = 16'hfe11;
#10;
address_ina = 74;
address_inb = 75;
data_ina = 16'hfd58;
data_inb = 16'h3f7;
#10;
address_ina = 76;
address_inb = 77;
data_ina = 16'h424;
data_inb = 16'hfccf;
#10;
address_ina = 78;
address_inb = 79;
data_ina = 16'h39c;
data_inb = 16'hfd59;
#10;
address_ina = 80;
address_inb = 81;
data_ina = 16'hff9f;
data_inb = 16'hfa2b;
#10;
address_ina = 82;
address_inb = 83;
data_ina = 16'h18c;
data_inb = 16'h20e;
#10;
address_ina = 84;
address_inb = 85;
data_ina = 16'h2bd;
data_inb = 16'h15;
#10;
address_ina = 86;
address_inb = 87;
data_ina = 16'hff9d;
data_inb = 16'h6c;
#10;
address_ina = 88;
address_inb = 89;
data_ina = 16'hfb22;
data_inb = 16'h1f7;
#10;
address_ina = 90;
address_inb = 91;
data_ina = 16'h55e;
data_inb = 16'h176;
#10;
address_ina = 92;
address_inb = 93;
data_ina = 16'h65c;
data_inb = 16'hfb17;
#10;
address_ina = 94;
address_inb = 95;
data_ina = 16'hfe6e;
data_inb = 16'h407;
#10;
address_ina = 96;
address_inb = 97;
data_ina = 16'hfb17;
data_inb = 16'hfd9f;
#10;
address_ina = 98;
address_inb = 99;
data_ina = 16'h61e;
data_inb = 16'hfb22;
#10;
address_ina = 100;
address_inb = 101;
data_ina = 16'h1e1;
data_inb = 16'h18f;
#10;
address_ina = 102;
address_inb = 103;
data_ina = 16'hfa29;
data_inb = 16'h3d1;
#10;
address_ina = 104;
address_inb = 105;
data_ina = 16'hfe15;
data_inb = 16'h65c;
#10;
address_ina = 106;
address_inb = 107;
data_ina = 16'h4ca;
data_inb = 16'hff60;
#10;
address_ina = 108;
address_inb = 109;
data_ina = 16'h486;
data_inb = 16'hff5b;
#10;
address_ina = 110;
address_inb = 111;
data_ina = 16'hfb1c;
data_inb = 16'h290;
#10;
address_ina = 112;
address_inb = 113;
data_ina = 16'hf9ea;
data_inb = 16'h205;
#10;
address_ina = 114;
address_inb = 115;
data_ina = 16'hfd6f;
data_inb = 16'h5d6;
#10;
address_ina = 116;
address_inb = 117;
data_ina = 16'hfb77;
data_inb = 16'hfca1;
#10;
address_ina = 118;
address_inb = 119;
data_ina = 16'hd6;
data_inb = 16'hffcb;
#10;
address_ina = 120;
address_inb = 121;
data_ina = 16'h55d;
data_inb = 16'hfae5;
#10;
address_ina = 122;
address_inb = 123;
data_ina = 16'hffc7;
data_inb = 16'hfdd7;
#10;
address_ina = 124;
address_inb = 125;
data_ina = 16'h144;
data_inb = 16'hfa9e;
#10;
address_ina = 126;
address_inb = 127;
data_ina = 16'hfab0;
data_inb = 16'h1ec;
#10;
address_ina = 128;
address_inb = 129;
data_ina = 16'hfdc7;
data_inb = 16'hfbfd;
#10;
address_ina = 130;
address_inb = 131;
data_ina = 16'hfbbf;
data_inb = 16'hff9a;
#10;
address_ina = 132;
address_inb = 133;
data_ina = 16'h66;
data_inb = 16'h3f6;
#10;
address_ina = 134;
address_inb = 135;
data_ina = 16'h2c9;
data_inb = 16'h198;
#10;
address_ina = 136;
address_inb = 137;
data_ina = 16'h51d;
data_inb = 16'h111;
#10;
address_ina = 138;
address_inb = 139;
data_ina = 16'hb3;
data_inb = 16'h32e;
#10;
address_ina = 140;
address_inb = 141;
data_ina = 16'h579;
data_inb = 16'hfc2a;
#10;
address_ina = 142;
address_inb = 143;
data_ina = 16'hfbbd;
data_inb = 16'hfcb2;
#10;
address_ina = 144;
address_inb = 145;
data_ina = 16'hfd0f;
data_inb = 16'hfc47;
#10;
address_ina = 146;
address_inb = 147;
data_ina = 16'hfc1d;
data_inb = 16'h1ad;
#10;
address_ina = 148;
address_inb = 149;
data_ina = 16'hff75;
data_inb = 16'hfa3c;
#10;
address_ina = 150;
address_inb = 151;
data_ina = 16'hfcd6;
data_inb = 16'h122;
#10;
address_ina = 152;
address_inb = 153;
data_ina = 16'hfa82;
data_inb = 16'h498;
#10;
address_ina = 154;
address_inb = 155;
data_ina = 16'hfbfb;
data_inb = 16'hfe16;
#10;
address_ina = 156;
address_inb = 157;
data_ina = 16'h91;
data_inb = 16'hfdcf;
#10;
address_ina = 158;
address_inb = 159;
data_ina = 16'hc7;
data_inb = 16'hf9ab;
#10;
address_ina = 160;
address_inb = 161;
data_ina = 16'hfea8;
data_inb = 16'hfc48;
#10;
address_ina = 162;
address_inb = 163;
data_ina = 16'hfa1f;
data_inb = 16'h393;
#10;
address_ina = 164;
address_inb = 165;
data_ina = 16'hfff2;
data_inb = 16'h27f;
#10;
address_ina = 166;
address_inb = 167;
data_ina = 16'h5a4;
data_inb = 16'h223;
#10;
address_ina = 168;
address_inb = 169;
data_ina = 16'hffb0;
data_inb = 16'h653;
#10;
address_ina = 170;
address_inb = 171;
data_ina = 16'hfe0c;
data_inb = 16'hfcf0;
#10;
address_ina = 172;
address_inb = 173;
data_ina = 16'h2a0;
data_inb = 16'hfd55;
#10;
address_ina = 174;
address_inb = 175;
data_ina = 16'hfd33;
data_inb = 16'h3fe;
#10;
address_ina = 176;
address_inb = 177;
data_ina = 16'h67a;
data_inb = 16'h608;
#10;
address_ina = 178;
address_inb = 179;
data_ina = 16'h1be;
data_inb = 16'hfd84;
#10;
address_ina = 180;
address_inb = 181;
data_ina = 16'hfb82;
data_inb = 16'h73;
#10;
address_ina = 182;
address_inb = 183;
data_ina = 16'h1f8;
data_inb = 16'h61c;
#10;
address_ina = 184;
address_inb = 185;
data_ina = 16'h472;
data_inb = 16'hfcd0;
#10;
address_ina = 186;
address_inb = 187;
data_ina = 16'h64b;
data_inb = 16'h3c7;
#10;
address_ina = 188;
address_inb = 189;
data_ina = 16'h5e7;
data_inb = 16'h2a7;
#10;
address_ina = 190;
address_inb = 191;
data_ina = 16'hfa35;
data_inb = 16'hff21;
#10;
address_ina = 192;
address_inb = 193;
data_ina = 16'hfee2;
data_inb = 16'h548;
#10;
address_ina = 194;
address_inb = 195;
data_ina = 16'h1e1;
data_inb = 16'h1cd;
#10;
address_ina = 196;
address_inb = 197;
data_ina = 16'hfeb8;
data_inb = 16'h425;
#10;
address_ina = 198;
address_inb = 199;
data_ina = 16'h143;
data_inb = 16'hfb96;
#10;
address_ina = 200;
address_inb = 201;
data_ina = 16'hfc71;
data_inb = 16'h1ed;
#10;
address_ina = 202;
address_inb = 203;
data_ina = 16'h4a9;
data_inb = 16'hfa43;
#10;
address_ina = 204;
address_inb = 205;
data_ina = 16'hffcc;
data_inb = 16'hfcb5;
#10;
address_ina = 206;
address_inb = 207;
data_ina = 16'hfc2b;
data_inb = 16'h10;
#10;
address_ina = 208;
address_inb = 209;
data_ina = 16'hfb95;
data_inb = 16'hfbe4;
#10;
address_ina = 210;
address_inb = 211;
data_ina = 16'hfc52;
data_inb = 16'hf9d9;
#10;
address_ina = 212;
address_inb = 213;
data_ina = 16'h1f0;
data_inb = 16'h5b9;
#10;
address_ina = 214;
address_inb = 215;
data_ina = 16'hfd46;
data_inb = 16'hfab5;
#10;
address_ina = 216;
address_inb = 217;
data_ina = 16'hfe48;
data_inb = 16'hf2;
#10;
address_ina = 218;
address_inb = 219;
data_ina = 16'h3f5;
data_inb = 16'hfa86;
#10;
address_ina = 220;
address_inb = 221;
data_ina = 16'hfad2;
data_inb = 16'hff14;
#10;
address_ina = 222;
address_inb = 223;
data_ina = 16'hee;
data_inb = 16'h2a8;
#10;
address_ina = 224;
address_inb = 225;
data_ina = 16'h561;
data_inb = 16'h45f;
#10;
address_ina = 226;
address_inb = 227;
data_ina = 16'h58b;
data_inb = 16'h64a;
#10;
address_ina = 228;
address_inb = 229;
data_ina = 16'h3eb;
data_inb = 16'hf9ea;
#10;
address_ina = 230;
address_inb = 231;
data_ina = 16'hfd93;
data_inb = 16'hfd61;
#10;
address_ina = 232;
address_inb = 233;
data_ina = 16'hfa18;
data_inb = 16'hfeff;
#10;
address_ina = 234;
address_inb = 235;
data_ina = 16'hfb1f;
data_inb = 16'h1cd;
#10;
address_ina = 236;
address_inb = 237;
data_ina = 16'hc7;
data_inb = 16'hfb81;
#10;
address_ina = 238;
address_inb = 239;
data_ina = 16'hf9c1;
data_inb = 16'h79;
#10;
address_ina = 240;
address_inb = 241;
data_ina = 16'h432;
data_inb = 16'hfbc6;
#10;
address_ina = 242;
address_inb = 243;
data_ina = 16'h5ea;
data_inb = 16'hfe43;
#10;
address_ina = 244;
address_inb = 245;
data_ina = 16'h517;
data_inb = 16'hf9f4;
#10;
address_ina = 246;
address_inb = 247;
data_ina = 16'h620;
data_inb = 16'hfbd3;
#10;
address_ina = 248;
address_inb = 249;
data_ina = 16'hfe0d;
data_inb = 16'hfec0;
#10;
address_ina = 250;
address_inb = 251;
data_ina = 16'hfb4b;
data_inb = 16'h497;
#10;
address_ina = 252;
address_inb = 253;
data_ina = 16'hfab9;
data_inb = 16'h239;
#10;
address_ina = 254;
address_inb = 255;
data_ina = 16'hff5f;
data_inb = 16'hfe69;
#10;
        wait(init_done);
        #30
        we = 0;
        // Start processing
         
		  #38000

        start = 0;



//        wait (wr_req);
//		  wait (!wr_req);
//		   rd_req = 1;
		  wait(done);
		  #20000
rd_req = 1;
        #70 
		  start = 1;
		 #80 
wait(rd_empty)
rd_req = 0;

$display("Finished the NTT test Number %d",test_num);
////Begin test number #76//////////////
rst = 1;

//#1000
start = 1;
mode = 1; //NTT 0 // INTT 1

// Reset for a few clock cycles

#1000

rst = 0;
test_num = test_num + 1;
#1000
we = 1;
address_ina = 0;
address_inb = 1;
data_ina = 16'hf9bc;
data_inb = 16'h28d;
#10;
address_ina = 2;
address_inb = 3;
data_ina = 16'hff92;
data_inb = 16'hf9ee;
#10;
address_ina = 4;
address_inb = 5;
data_ina = 16'h36;
data_inb = 16'hfef9;
#10;
address_ina = 6;
address_inb = 7;
data_ina = 16'hfbf0;
data_inb = 16'hf9dc;
#10;
address_ina = 8;
address_inb = 9;
data_ina = 16'hae;
data_inb = 16'hfed5;
#10;
address_ina = 10;
address_inb = 11;
data_ina = 16'h5fb;
data_inb = 16'hfe2e;
#10;
address_ina = 12;
address_inb = 13;
data_ina = 16'hf5;
data_inb = 16'hfa89;
#10;
address_ina = 14;
address_inb = 15;
data_ina = 16'hfc3d;
data_inb = 16'h129;
#10;
address_ina = 16;
address_inb = 17;
data_ina = 16'hfc8f;
data_inb = 16'hfce4;
#10;
address_ina = 18;
address_inb = 19;
data_ina = 16'h1e7;
data_inb = 16'h540;
#10;
address_ina = 20;
address_inb = 21;
data_ina = 16'hfa29;
data_inb = 16'h61e;
#10;
address_ina = 22;
address_inb = 23;
data_ina = 16'h4;
data_inb = 16'hfced;
#10;
address_ina = 24;
address_inb = 25;
data_ina = 16'hfd9b;
data_inb = 16'hfa8b;
#10;
address_ina = 26;
address_inb = 27;
data_ina = 16'h1dd;
data_inb = 16'hfce6;
#10;
address_ina = 28;
address_inb = 29;
data_ina = 16'h301;
data_inb = 16'h1d3;
#10;
address_ina = 30;
address_inb = 31;
data_ina = 16'h2bc;
data_inb = 16'hff53;
#10;
address_ina = 32;
address_inb = 33;
data_ina = 16'h584;
data_inb = 16'h27b;
#10;
address_ina = 34;
address_inb = 35;
data_ina = 16'h31e;
data_inb = 16'hfc1c;
#10;
address_ina = 36;
address_inb = 37;
data_ina = 16'hff07;
data_inb = 16'h4a5;
#10;
address_ina = 38;
address_inb = 39;
data_ina = 16'hfd03;
data_inb = 16'h500;
#10;
address_ina = 40;
address_inb = 41;
data_ina = 16'hfb84;
data_inb = 16'h383;
#10;
address_ina = 42;
address_inb = 43;
data_ina = 16'hfe9a;
data_inb = 16'hfa5d;
#10;
address_ina = 44;
address_inb = 45;
data_ina = 16'h1ed;
data_inb = 16'h2d5;
#10;
address_ina = 46;
address_inb = 47;
data_ina = 16'h218;
data_inb = 16'h228;
#10;
address_ina = 48;
address_inb = 49;
data_ina = 16'h156;
data_inb = 16'hfacf;
#10;
address_ina = 50;
address_inb = 51;
data_ina = 16'hfe22;
data_inb = 16'hfb6b;
#10;
address_ina = 52;
address_inb = 53;
data_ina = 16'h206;
data_inb = 16'hfe4e;
#10;
address_ina = 54;
address_inb = 55;
data_ina = 16'hfdbe;
data_inb = 16'h1ff;
#10;
address_ina = 56;
address_inb = 57;
data_ina = 16'h221;
data_inb = 16'h2be;
#10;
address_ina = 58;
address_inb = 59;
data_ina = 16'h2fa;
data_inb = 16'h63;
#10;
address_ina = 60;
address_inb = 61;
data_ina = 16'hfb2a;
data_inb = 16'hfe3a;
#10;
address_ina = 62;
address_inb = 63;
data_ina = 16'hfe41;
data_inb = 16'hff98;
#10;
address_ina = 64;
address_inb = 65;
data_ina = 16'h599;
data_inb = 16'hffa8;
#10;
address_ina = 66;
address_inb = 67;
data_ina = 16'hfe83;
data_inb = 16'hff0e;
#10;
address_ina = 68;
address_inb = 69;
data_ina = 16'h4f4;
data_inb = 16'h5d0;
#10;
address_ina = 70;
address_inb = 71;
data_ina = 16'hfbe6;
data_inb = 16'h146;
#10;
address_ina = 72;
address_inb = 73;
data_ina = 16'h635;
data_inb = 16'h4ae;
#10;
address_ina = 74;
address_inb = 75;
data_ina = 16'hf9d6;
data_inb = 16'h8d;
#10;
address_ina = 76;
address_inb = 77;
data_ina = 16'hfae6;
data_inb = 16'h1b;
#10;
address_ina = 78;
address_inb = 79;
data_ina = 16'hfd9b;
data_inb = 16'hfa63;
#10;
address_ina = 80;
address_inb = 81;
data_ina = 16'hff41;
data_inb = 16'hfa1d;
#10;
address_ina = 82;
address_inb = 83;
data_ina = 16'hfdcc;
data_inb = 16'h2d;
#10;
address_ina = 84;
address_inb = 85;
data_ina = 16'h534;
data_inb = 16'h201;
#10;
address_ina = 86;
address_inb = 87;
data_ina = 16'hfc;
data_inb = 16'h151;
#10;
address_ina = 88;
address_inb = 89;
data_ina = 16'h471;
data_inb = 16'h67;
#10;
address_ina = 90;
address_inb = 91;
data_ina = 16'h369;
data_inb = 16'h59d;
#10;
address_ina = 92;
address_inb = 93;
data_ina = 16'hfd47;
data_inb = 16'h2ea;
#10;
address_ina = 94;
address_inb = 95;
data_ina = 16'hffde;
data_inb = 16'h420;
#10;
address_ina = 96;
address_inb = 97;
data_ina = 16'h592;
data_inb = 16'hff80;
#10;
address_ina = 98;
address_inb = 99;
data_ina = 16'hfb5b;
data_inb = 16'h65;
#10;
address_ina = 100;
address_inb = 101;
data_ina = 16'hfcab;
data_inb = 16'hfc7f;
#10;
address_ina = 102;
address_inb = 103;
data_ina = 16'h49;
data_inb = 16'hfbe3;
#10;
address_ina = 104;
address_inb = 105;
data_ina = 16'hfb82;
data_inb = 16'hfe6e;
#10;
address_ina = 106;
address_inb = 107;
data_ina = 16'h1ce;
data_inb = 16'h286;
#10;
address_ina = 108;
address_inb = 109;
data_ina = 16'h93;
data_inb = 16'h4cc;
#10;
address_ina = 110;
address_inb = 111;
data_ina = 16'hffb0;
data_inb = 16'h596;
#10;
address_ina = 112;
address_inb = 113;
data_ina = 16'h385;
data_inb = 16'h505;
#10;
address_ina = 114;
address_inb = 115;
data_ina = 16'h357;
data_inb = 16'h39a;
#10;
address_ina = 116;
address_inb = 117;
data_ina = 16'hff6e;
data_inb = 16'h364;
#10;
address_ina = 118;
address_inb = 119;
data_ina = 16'hffcc;
data_inb = 16'hfc2f;
#10;
address_ina = 120;
address_inb = 121;
data_ina = 16'h48;
data_inb = 16'h227;
#10;
address_ina = 122;
address_inb = 123;
data_ina = 16'hfc99;
data_inb = 16'h488;
#10;
address_ina = 124;
address_inb = 125;
data_ina = 16'h2ac;
data_inb = 16'hfc31;
#10;
address_ina = 126;
address_inb = 127;
data_ina = 16'hfbf4;
data_inb = 16'hfcbe;
#10;
address_ina = 128;
address_inb = 129;
data_ina = 16'hfa00;
data_inb = 16'hfdcf;
#10;
address_ina = 130;
address_inb = 131;
data_ina = 16'hdd;
data_inb = 16'h35d;
#10;
address_ina = 132;
address_inb = 133;
data_ina = 16'hfb8d;
data_inb = 16'hfdd6;
#10;
address_ina = 134;
address_inb = 135;
data_ina = 16'h3e4;
data_inb = 16'hf9e7;
#10;
address_ina = 136;
address_inb = 137;
data_ina = 16'hfbbc;
data_inb = 16'h442;
#10;
address_ina = 138;
address_inb = 139;
data_ina = 16'h45d;
data_inb = 16'hfa18;
#10;
address_ina = 140;
address_inb = 141;
data_ina = 16'h136;
data_inb = 16'hfaab;
#10;
address_ina = 142;
address_inb = 143;
data_ina = 16'hfd99;
data_inb = 16'hff28;
#10;
address_ina = 144;
address_inb = 145;
data_ina = 16'hfdb5;
data_inb = 16'hfabb;
#10;
address_ina = 146;
address_inb = 147;
data_ina = 16'hfa90;
data_inb = 16'h7;
#10;
address_ina = 148;
address_inb = 149;
data_ina = 16'h1b8;
data_inb = 16'h8a;
#10;
address_ina = 150;
address_inb = 151;
data_ina = 16'hfbeb;
data_inb = 16'hff53;
#10;
address_ina = 152;
address_inb = 153;
data_ina = 16'h17b;
data_inb = 16'hfef8;
#10;
address_ina = 154;
address_inb = 155;
data_ina = 16'h51b;
data_inb = 16'hffd8;
#10;
address_ina = 156;
address_inb = 157;
data_ina = 16'hfbc9;
data_inb = 16'h2c0;
#10;
address_ina = 158;
address_inb = 159;
data_ina = 16'h102;
data_inb = 16'h545;
#10;
address_ina = 160;
address_inb = 161;
data_ina = 16'h328;
data_inb = 16'hf9ae;
#10;
address_ina = 162;
address_inb = 163;
data_ina = 16'hfe55;
data_inb = 16'hfca4;
#10;
address_ina = 164;
address_inb = 165;
data_ina = 16'hfef3;
data_inb = 16'h517;
#10;
address_ina = 166;
address_inb = 167;
data_ina = 16'h395;
data_inb = 16'hfe38;
#10;
address_ina = 168;
address_inb = 169;
data_ina = 16'h444;
data_inb = 16'hff80;
#10;
address_ina = 170;
address_inb = 171;
data_ina = 16'hfff6;
data_inb = 16'h116;
#10;
address_ina = 172;
address_inb = 173;
data_ina = 16'h400;
data_inb = 16'hf996;
#10;
address_ina = 174;
address_inb = 175;
data_ina = 16'hff6f;
data_inb = 16'hfeed;
#10;
address_ina = 176;
address_inb = 177;
data_ina = 16'h3f7;
data_inb = 16'hfc94;
#10;
address_ina = 178;
address_inb = 179;
data_ina = 16'h4e;
data_inb = 16'hf9c7;
#10;
address_ina = 180;
address_inb = 181;
data_ina = 16'hae;
data_inb = 16'h5f8;
#10;
address_ina = 182;
address_inb = 183;
data_ina = 16'hfeb5;
data_inb = 16'hfc2b;
#10;
address_ina = 184;
address_inb = 185;
data_ina = 16'hff6a;
data_inb = 16'h3b3;
#10;
address_ina = 186;
address_inb = 187;
data_ina = 16'hfee4;
data_inb = 16'hffb8;
#10;
address_ina = 188;
address_inb = 189;
data_ina = 16'h238;
data_inb = 16'hfa37;
#10;
address_ina = 190;
address_inb = 191;
data_ina = 16'h305;
data_inb = 16'hfb57;
#10;
address_ina = 192;
address_inb = 193;
data_ina = 16'hfae4;
data_inb = 16'hfd8f;
#10;
address_ina = 194;
address_inb = 195;
data_ina = 16'hfe2c;
data_inb = 16'h17b;
#10;
address_ina = 196;
address_inb = 197;
data_ina = 16'hfc41;
data_inb = 16'hfa93;
#10;
address_ina = 198;
address_inb = 199;
data_ina = 16'h42;
data_inb = 16'h58e;
#10;
address_ina = 200;
address_inb = 201;
data_ina = 16'hfe09;
data_inb = 16'hff17;
#10;
address_ina = 202;
address_inb = 203;
data_ina = 16'h566;
data_inb = 16'h669;
#10;
address_ina = 204;
address_inb = 205;
data_ina = 16'hfe6b;
data_inb = 16'hf9d2;
#10;
address_ina = 206;
address_inb = 207;
data_ina = 16'h2c8;
data_inb = 16'hfd0e;
#10;
address_ina = 208;
address_inb = 209;
data_ina = 16'hf3;
data_inb = 16'hfc9c;
#10;
address_ina = 210;
address_inb = 211;
data_ina = 16'h489;
data_inb = 16'hfa7b;
#10;
address_ina = 212;
address_inb = 213;
data_ina = 16'hfe3f;
data_inb = 16'h4e7;
#10;
address_ina = 214;
address_inb = 215;
data_ina = 16'h3e;
data_inb = 16'hfcb6;
#10;
address_ina = 216;
address_inb = 217;
data_ina = 16'hfb42;
data_inb = 16'hfa01;
#10;
address_ina = 218;
address_inb = 219;
data_ina = 16'hfd51;
data_inb = 16'h2d9;
#10;
address_ina = 220;
address_inb = 221;
data_ina = 16'hfd37;
data_inb = 16'h48e;
#10;
address_ina = 222;
address_inb = 223;
data_ina = 16'h5a2;
data_inb = 16'hfcda;
#10;
address_ina = 224;
address_inb = 225;
data_ina = 16'hfd1d;
data_inb = 16'h173;
#10;
address_ina = 226;
address_inb = 227;
data_ina = 16'hff9d;
data_inb = 16'h536;
#10;
address_ina = 228;
address_inb = 229;
data_ina = 16'hfcf6;
data_inb = 16'h568;
#10;
address_ina = 230;
address_inb = 231;
data_ina = 16'hfe50;
data_inb = 16'hfb10;
#10;
address_ina = 232;
address_inb = 233;
data_ina = 16'hfd34;
data_inb = 16'hfc69;
#10;
address_ina = 234;
address_inb = 235;
data_ina = 16'h467;
data_inb = 16'h554;
#10;
address_ina = 236;
address_inb = 237;
data_ina = 16'h47c;
data_inb = 16'hfcfc;
#10;
address_ina = 238;
address_inb = 239;
data_ina = 16'hfa89;
data_inb = 16'hfbb4;
#10;
address_ina = 240;
address_inb = 241;
data_ina = 16'hff68;
data_inb = 16'h2b5;
#10;
address_ina = 242;
address_inb = 243;
data_ina = 16'hfcbd;
data_inb = 16'hfb07;
#10;
address_ina = 244;
address_inb = 245;
data_ina = 16'h446;
data_inb = 16'h3de;
#10;
address_ina = 246;
address_inb = 247;
data_ina = 16'hff38;
data_inb = 16'hfb3b;
#10;
address_ina = 248;
address_inb = 249;
data_ina = 16'hfab7;
data_inb = 16'hfaa3;
#10;
address_ina = 250;
address_inb = 251;
data_ina = 16'hff5e;
data_inb = 16'h4f9;
#10;
address_ina = 252;
address_inb = 253;
data_ina = 16'hf9ae;
data_inb = 16'h2f8;
#10;
address_ina = 254;
address_inb = 255;
data_ina = 16'h3a9;
data_inb = 16'h633;
#10;
        wait(init_done);
        #30
        we = 0;
        // Start processing
         
		  #38000

        start = 0;



//        wait (wr_req);
//		  wait (!wr_req);
//		   rd_req = 1;
		  wait(done);
		  #20000
rd_req = 1;
        #70 
		  start = 1;
		 #80 
wait(rd_empty)
rd_req = 0;

$display("Finished the NTT test Number %d",test_num);
////Begin test number #77//////////////
rst = 1;

//#1000
start = 1;
mode = 0; //NTT 0 // INTT 1

// Reset for a few clock cycles

#1000

rst = 0;
test_num = test_num + 1;
#1000
we = 1;
address_ina = 0;
address_inb = 1;
data_ina = 16'h979;
data_inb = 16'hc8c;
#10;
address_ina = 2;
address_inb = 3;
data_ina = 16'hda;
data_inb = 16'h754;
#10;
address_ina = 4;
address_inb = 5;
data_ina = 16'h938;
data_inb = 16'h74a;
#10;
address_ina = 6;
address_inb = 7;
data_ina = 16'h499;
data_inb = 16'ha94;
#10;
address_ina = 8;
address_inb = 9;
data_ina = 16'h30c;
data_inb = 16'h5f1;
#10;
address_ina = 10;
address_inb = 11;
data_ina = 16'hcc0;
data_inb = 16'hb8b;
#10;
address_ina = 12;
address_inb = 13;
data_ina = 16'hc00;
data_inb = 16'h5e;
#10;
address_ina = 14;
address_inb = 15;
data_ina = 16'h5aa;
data_inb = 16'h6df;
#10;
address_ina = 16;
address_inb = 17;
data_ina = 16'h215;
data_inb = 16'h62c;
#10;
address_ina = 18;
address_inb = 19;
data_ina = 16'h66a;
data_inb = 16'h243;
#10;
address_ina = 20;
address_inb = 21;
data_ina = 16'h8ea;
data_inb = 16'ha05;
#10;
address_ina = 22;
address_inb = 23;
data_ina = 16'h208;
data_inb = 16'hc3;
#10;
address_ina = 24;
address_inb = 25;
data_ina = 16'h57c;
data_inb = 16'h962;
#10;
address_ina = 26;
address_inb = 27;
data_ina = 16'h159;
data_inb = 16'hd3;
#10;
address_ina = 28;
address_inb = 29;
data_ina = 16'ha77;
data_inb = 16'h76b;
#10;
address_ina = 30;
address_inb = 31;
data_ina = 16'h17;
data_inb = 16'h86b;
#10;
address_ina = 32;
address_inb = 33;
data_ina = 16'hc4e;
data_inb = 16'hc37;
#10;
address_ina = 34;
address_inb = 35;
data_ina = 16'h9ce;
data_inb = 16'h6df;
#10;
address_ina = 36;
address_inb = 37;
data_ina = 16'h821;
data_inb = 16'hba5;
#10;
address_ina = 38;
address_inb = 39;
data_ina = 16'hcf1;
data_inb = 16'h7;
#10;
address_ina = 40;
address_inb = 41;
data_ina = 16'h33d;
data_inb = 16'h6e2;
#10;
address_ina = 42;
address_inb = 43;
data_ina = 16'h596;
data_inb = 16'h246;
#10;
address_ina = 44;
address_inb = 45;
data_ina = 16'h2a7;
data_inb = 16'h6bb;
#10;
address_ina = 46;
address_inb = 47;
data_ina = 16'h4ea;
data_inb = 16'h55c;
#10;
address_ina = 48;
address_inb = 49;
data_ina = 16'h925;
data_inb = 16'h22f;
#10;
address_ina = 50;
address_inb = 51;
data_ina = 16'h966;
data_inb = 16'h3f0;
#10;
address_ina = 52;
address_inb = 53;
data_ina = 16'h22c;
data_inb = 16'h2e5;
#10;
address_ina = 54;
address_inb = 55;
data_ina = 16'h583;
data_inb = 16'h962;
#10;
address_ina = 56;
address_inb = 57;
data_ina = 16'h851;
data_inb = 16'h96c;
#10;
address_ina = 58;
address_inb = 59;
data_ina = 16'h1a3;
data_inb = 16'h1c1;
#10;
address_ina = 60;
address_inb = 61;
data_ina = 16'h9d4;
data_inb = 16'h878;
#10;
address_ina = 62;
address_inb = 63;
data_ina = 16'h239;
data_inb = 16'hb16;
#10;
address_ina = 64;
address_inb = 65;
data_ina = 16'haef;
data_inb = 16'h8b0;
#10;
address_ina = 66;
address_inb = 67;
data_ina = 16'hb92;
data_inb = 16'hba8;
#10;
address_ina = 68;
address_inb = 69;
data_ina = 16'h945;
data_inb = 16'h3a2;
#10;
address_ina = 70;
address_inb = 71;
data_ina = 16'h650;
data_inb = 16'h785;
#10;
address_ina = 72;
address_inb = 73;
data_ina = 16'h8d3;
data_inb = 16'h91b;
#10;
address_ina = 74;
address_inb = 75;
data_ina = 16'h496;
data_inb = 16'h8d3;
#10;
address_ina = 76;
address_inb = 77;
data_ina = 16'h378;
data_inb = 16'hcc3;
#10;
address_ina = 78;
address_inb = 79;
data_ina = 16'h3d9;
data_inb = 16'h63c;
#10;
address_ina = 80;
address_inb = 81;
data_ina = 16'hb06;
data_inb = 16'h7b5;
#10;
address_ina = 82;
address_inb = 83;
data_ina = 16'h458;
data_inb = 16'h7fd;
#10;
address_ina = 84;
address_inb = 85;
data_ina = 16'hbe3;
data_inb = 16'h6b;
#10;
address_ina = 86;
address_inb = 87;
data_ina = 16'hb54;
data_inb = 16'h1d;
#10;
address_ina = 88;
address_inb = 89;
data_ina = 16'h183;
data_inb = 16'h612;
#10;
address_ina = 90;
address_inb = 91;
data_ina = 16'h22c;
data_inb = 16'h10b;
#10;
address_ina = 92;
address_inb = 93;
data_ina = 16'h5e;
data_inb = 16'h58;
#10;
address_ina = 94;
address_inb = 95;
data_ina = 16'h72d;
data_inb = 16'haa1;
#10;
address_ina = 96;
address_inb = 97;
data_ina = 16'h9e1;
data_inb = 16'h9f;
#10;
address_ina = 98;
address_inb = 99;
data_ina = 16'ha40;
data_inb = 16'hb3d;
#10;
address_ina = 100;
address_inb = 101;
data_ina = 16'hb9;
data_inb = 16'h7f3;
#10;
address_ina = 102;
address_inb = 103;
data_ina = 16'h354;
data_inb = 16'ha70;
#10;
address_ina = 104;
address_inb = 105;
data_ina = 16'ha40;
data_inb = 16'h7b9;
#10;
address_ina = 106;
address_inb = 107;
data_ina = 16'h7f;
data_inb = 16'h9bd;
#10;
address_ina = 108;
address_inb = 109;
data_ina = 16'hbd3;
data_inb = 16'hb67;
#10;
address_ina = 110;
address_inb = 111;
data_ina = 16'h7f;
data_inb = 16'h9c7;
#10;
address_ina = 112;
address_inb = 113;
data_ina = 16'h344;
data_inb = 16'h101;
#10;
address_ina = 114;
address_inb = 115;
data_ina = 16'h91b;
data_inb = 16'h96f;
#10;
address_ina = 116;
address_inb = 117;
data_ina = 16'h580;
data_inb = 16'h740;
#10;
address_ina = 118;
address_inb = 119;
data_ina = 16'h7d6;
data_inb = 16'h8ed;
#10;
address_ina = 120;
address_inb = 121;
data_ina = 16'h831;
data_inb = 16'hce7;
#10;
address_ina = 122;
address_inb = 123;
data_ina = 16'h16c;
data_inb = 16'ha0c;
#10;
address_ina = 124;
address_inb = 125;
data_ina = 16'ha3;
data_inb = 16'h2b8;
#10;
address_ina = 126;
address_inb = 127;
data_ina = 16'h966;
data_inb = 16'h250;
#10;
address_ina = 128;
address_inb = 129;
data_ina = 16'h319;
data_inb = 16'h55;
#10;
address_ina = 130;
address_inb = 131;
data_ina = 16'hc75;
data_inb = 16'h632;
#10;
address_ina = 132;
address_inb = 133;
data_ina = 16'h4d7;
data_inb = 16'ha15;
#10;
address_ina = 134;
address_inb = 135;
data_ina = 16'h9f2;
data_inb = 16'h1f8;
#10;
address_ina = 136;
address_inb = 137;
data_ina = 16'h78e;
data_inb = 16'h656;
#10;
address_ina = 138;
address_inb = 139;
data_ina = 16'h3b;
data_inb = 16'h925;
#10;
address_ina = 140;
address_inb = 141;
data_ina = 16'h2db;
data_inb = 16'hb6;
#10;
address_ina = 142;
address_inb = 143;
data_ina = 16'h559;
data_inb = 16'h6c5;
#10;
address_ina = 144;
address_inb = 145;
data_ina = 16'h6f9;
data_inb = 16'h256;
#10;
address_ina = 146;
address_inb = 147;
data_ina = 16'hcc6;
data_inb = 16'hb0;
#10;
address_ina = 148;
address_inb = 149;
data_ina = 16'ha02;
data_inb = 16'h104;
#10;
address_ina = 150;
address_inb = 151;
data_ina = 16'h458;
data_inb = 16'h3e9;
#10;
address_ina = 152;
address_inb = 153;
data_ina = 16'h9ff;
data_inb = 16'h7b9;
#10;
address_ina = 154;
address_inb = 155;
data_ina = 16'hea;
data_inb = 16'h6ae;
#10;
address_ina = 156;
address_inb = 157;
data_ina = 16'h9b7;
data_inb = 16'h34a;
#10;
address_ina = 158;
address_inb = 159;
data_ina = 16'h64c;
data_inb = 16'h3e;
#10;
address_ina = 160;
address_inb = 161;
data_ina = 16'h703;
data_inb = 16'hced;
#10;
address_ina = 162;
address_inb = 163;
data_ina = 16'h125;
data_inb = 16'h9c1;
#10;
address_ina = 164;
address_inb = 165;
data_ina = 16'h78b;
data_inb = 16'hb67;
#10;
address_ina = 166;
address_inb = 167;
data_ina = 16'h3b;
data_inb = 16'h183;
#10;
address_ina = 168;
address_inb = 169;
data_ina = 16'hca3;
data_inb = 16'h8b3;
#10;
address_ina = 170;
address_inb = 171;
data_ina = 16'h602;
data_inb = 16'hb6;
#10;
address_ina = 172;
address_inb = 173;
data_ina = 16'h9a0;
data_inb = 16'h68;
#10;
address_ina = 174;
address_inb = 175;
data_ina = 16'h246;
data_inb = 16'h788;
#10;
address_ina = 176;
address_inb = 177;
data_ina = 16'hbf6;
data_inb = 16'h99a;
#10;
address_ina = 178;
address_inb = 179;
data_ina = 16'h7c9;
data_inb = 16'h9e8;
#10;
address_ina = 180;
address_inb = 181;
data_ina = 16'hced;
data_inb = 16'h858;
#10;
address_ina = 182;
address_inb = 183;
data_ina = 16'h67d;
data_inb = 16'h173;
#10;
address_ina = 184;
address_inb = 185;
data_ina = 16'h79f;
data_inb = 16'h132;
#10;
address_ina = 186;
address_inb = 187;
data_ina = 16'h55c;
data_inb = 16'h559;
#10;
address_ina = 188;
address_inb = 189;
data_ina = 16'h525;
data_inb = 16'h17;
#10;
address_ina = 190;
address_inb = 191;
data_ina = 16'h545;
data_inb = 16'h385;
#10;
address_ina = 192;
address_inb = 193;
data_ina = 16'hbdc;
data_inb = 16'h737;
#10;
address_ina = 194;
address_inb = 195;
data_ina = 16'h3e0;
data_inb = 16'h778;
#10;
address_ina = 196;
address_inb = 197;
data_ina = 16'h38e;
data_inb = 16'h868;
#10;
address_ina = 198;
address_inb = 199;
data_ina = 16'h417;
data_inb = 16'hc10;
#10;
address_ina = 200;
address_inb = 201;
data_ina = 16'h706;
data_inb = 16'h114;
#10;
address_ina = 202;
address_inb = 203;
data_ina = 16'h294;
data_inb = 16'h12b;
#10;
address_ina = 204;
address_inb = 205;
data_ina = 16'h4e4;
data_inb = 16'h53b;
#10;
address_ina = 206;
address_inb = 207;
data_ina = 16'h583;
data_inb = 16'h3e;
#10;
address_ina = 208;
address_inb = 209;
data_ina = 16'hb23;
data_inb = 16'h3;
#10;
address_ina = 210;
address_inb = 211;
data_ina = 16'hcc3;
data_inb = 16'h417;
#10;
address_ina = 212;
address_inb = 213;
data_ina = 16'h5c7;
data_inb = 16'h99;
#10;
address_ina = 214;
address_inb = 215;
data_ina = 16'hb95;
data_inb = 16'h2df;
#10;
address_ina = 216;
address_inb = 217;
data_ina = 16'h76e;
data_inb = 16'hacf;
#10;
address_ina = 218;
address_inb = 219;
data_ina = 16'h3bf;
data_inb = 16'h7c9;
#10;
address_ina = 220;
address_inb = 221;
data_ina = 16'h993;
data_inb = 16'hcfa;
#10;
address_ina = 222;
address_inb = 223;
data_ina = 16'h27d;
data_inb = 16'h89c;
#10;
address_ina = 224;
address_inb = 225;
data_ina = 16'h82e;
data_inb = 16'h38e;
#10;
address_ina = 226;
address_inb = 227;
data_ina = 16'h395;
data_inb = 16'h36b;
#10;
address_ina = 228;
address_inb = 229;
data_ina = 16'hb5e;
data_inb = 16'h9e1;
#10;
address_ina = 230;
address_inb = 231;
data_ina = 16'hcf1;
data_inb = 16'h249;
#10;
address_ina = 232;
address_inb = 233;
data_ina = 16'h87c;
data_inb = 16'hbcf;
#10;
address_ina = 234;
address_inb = 235;
data_ina = 16'h5d7;
data_inb = 16'h17c;
#10;
address_ina = 236;
address_inb = 237;
data_ina = 16'h39f;
data_inb = 16'h7ac;
#10;
address_ina = 238;
address_inb = 239;
data_ina = 16'h875;
data_inb = 16'hd7;
#10;
address_ina = 240;
address_inb = 241;
data_ina = 16'h128;
data_inb = 16'hcb0;
#10;
address_ina = 242;
address_inb = 243;
data_ina = 16'hc9c;
data_inb = 16'hb09;
#10;
address_ina = 244;
address_inb = 245;
data_ina = 16'h6c2;
data_inb = 16'h7b5;
#10;
address_ina = 246;
address_inb = 247;
data_ina = 16'hc92;
data_inb = 16'hbd6;
#10;
address_ina = 248;
address_inb = 249;
data_ina = 16'h5ca;
data_inb = 16'ha19;
#10;
address_ina = 250;
address_inb = 251;
data_ina = 16'h35e;
data_inb = 16'h319;
#10;
address_ina = 252;
address_inb = 253;
data_ina = 16'hf4;
data_inb = 16'h872;
#10;
address_ina = 254;
address_inb = 255;
data_ina = 16'h2e8;
data_inb = 16'h5a0;
#10;
        wait(init_done);
        #30
        we = 0;
        // Start processing
         
		  #38000

        start = 0;



//        wait (wr_req);
//		  wait (!wr_req);
//		   rd_req = 1;
		  wait(done);
		  #20000
rd_req = 1;
        #70 
		  start = 1;
		 #80 
wait(rd_empty)
rd_req = 0;

$display("Finished the NTT test Number %d",test_num);
////Begin test number #78//////////////
rst = 1;

//#1000
start = 1;
mode = 0; //NTT 0 // INTT 1

// Reset for a few clock cycles

#1000

rst = 0;
test_num = test_num + 1;
#1000
we = 1;
address_ina = 0;
address_inb = 1;
data_ina = 16'h25d;
data_inb = 16'hfa;
#10;
address_ina = 2;
address_inb = 3;
data_ina = 16'h1c1;
data_inb = 16'hc1d;
#10;
address_ina = 4;
address_inb = 5;
data_ina = 16'hca;
data_inb = 16'h34;
#10;
address_ina = 6;
address_inb = 7;
data_ina = 16'h58;
data_inb = 16'h85;
#10;
address_ina = 8;
address_inb = 9;
data_ina = 16'h6d2;
data_inb = 16'hc1d;
#10;
address_ina = 10;
address_inb = 11;
data_ina = 16'h1a3;
data_inb = 16'h5b0;
#10;
address_ina = 12;
address_inb = 13;
data_ina = 16'h38b;
data_inb = 16'h2ec;
#10;
address_ina = 14;
address_inb = 15;
data_ina = 16'hb98;
data_inb = 16'hd3;
#10;
address_ina = 16;
address_inb = 17;
data_ina = 16'h1ce;
data_inb = 16'h807;
#10;
address_ina = 18;
address_inb = 19;
data_ina = 16'h807;
data_inb = 16'h81d;
#10;
address_ina = 20;
address_inb = 21;
data_ina = 16'h885;
data_inb = 16'h7f6;
#10;
address_ina = 22;
address_inb = 23;
data_ina = 16'h555;
data_inb = 16'h208;
#10;
address_ina = 24;
address_inb = 25;
data_ina = 16'h81a;
data_inb = 16'h489;
#10;
address_ina = 26;
address_inb = 27;
data_ina = 16'ha2c;
data_inb = 16'h20b;
#10;
address_ina = 28;
address_inb = 29;
data_ina = 16'h593;
data_inb = 16'hc10;
#10;
address_ina = 30;
address_inb = 31;
data_ina = 16'h4d0;
data_inb = 16'hc2a;
#10;
address_ina = 32;
address_inb = 33;
data_ina = 16'h367;
data_inb = 16'h51e;
#10;
address_ina = 34;
address_inb = 35;
data_ina = 16'h9e8;
data_inb = 16'h7e0;
#10;
address_ina = 36;
address_inb = 37;
data_ina = 16'h35e;
data_inb = 16'habb;
#10;
address_ina = 38;
address_inb = 39;
data_ina = 16'h5c4;
data_inb = 16'h225;
#10;
address_ina = 40;
address_inb = 41;
data_ina = 16'h751;
data_inb = 16'hb71;
#10;
address_ina = 42;
address_inb = 43;
data_ina = 16'hac2;
data_inb = 16'h7d3;
#10;
address_ina = 44;
address_inb = 45;
data_ina = 16'h4cd;
data_inb = 16'h6dc;
#10;
address_ina = 46;
address_inb = 47;
data_ina = 16'h4ca;
data_inb = 16'h11e;
#10;
address_ina = 48;
address_inb = 49;
data_ina = 16'h83e;
data_inb = 16'h882;
#10;
address_ina = 50;
address_inb = 51;
data_ina = 16'h5e1;
data_inb = 16'h5ba;
#10;
address_ina = 52;
address_inb = 53;
data_ina = 16'h925;
data_inb = 16'h821;
#10;
address_ina = 54;
address_inb = 55;
data_ina = 16'h511;
data_inb = 16'h266;
#10;
address_ina = 56;
address_inb = 57;
data_ina = 16'h945;
data_inb = 16'h2b4;
#10;
address_ina = 58;
address_inb = 59;
data_ina = 16'h9d1;
data_inb = 16'h37e;
#10;
address_ina = 60;
address_inb = 61;
data_ina = 16'h709;
data_inb = 16'h507;
#10;
address_ina = 62;
address_inb = 63;
data_ina = 16'h95c;
data_inb = 16'h316;
#10;
address_ina = 64;
address_inb = 65;
data_ina = 16'h320;
data_inb = 16'h8ea;
#10;
address_ina = 66;
address_inb = 67;
data_ina = 16'h43b;
data_inb = 16'hcb6;
#10;
address_ina = 68;
address_inb = 69;
data_ina = 16'h9b0;
data_inb = 16'h7ac;
#10;
address_ina = 70;
address_inb = 71;
data_ina = 16'hb10;
data_inb = 16'h4ca;
#10;
address_ina = 72;
address_inb = 73;
data_ina = 16'hce7;
data_inb = 16'h434;
#10;
address_ina = 74;
address_inb = 75;
data_ina = 16'ha08;
data_inb = 16'ha91;
#10;
address_ina = 76;
address_inb = 77;
data_ina = 16'h3d6;
data_inb = 16'h11e;
#10;
address_ina = 78;
address_inb = 79;
data_ina = 16'h186;
data_inb = 16'ha77;
#10;
address_ina = 80;
address_inb = 81;
data_ina = 16'h138;
data_inb = 16'hc6b;
#10;
address_ina = 82;
address_inb = 83;
data_ina = 16'hea;
data_inb = 16'hf4;
#10;
address_ina = 84;
address_inb = 85;
data_ina = 16'h496;
data_inb = 16'hb5e;
#10;
address_ina = 86;
address_inb = 87;
data_ina = 16'h2fc;
data_inb = 16'h88c;
#10;
address_ina = 88;
address_inb = 89;
data_ina = 16'h41a;
data_inb = 16'hbfd;
#10;
address_ina = 90;
address_inb = 91;
data_ina = 16'h605;
data_inb = 16'h7d6;
#10;
address_ina = 92;
address_inb = 93;
data_ina = 16'h47c;
data_inb = 16'h7;
#10;
address_ina = 94;
address_inb = 95;
data_ina = 16'hc2a;
data_inb = 16'h896;
#10;
address_ina = 96;
address_inb = 97;
data_ina = 16'h4bd;
data_inb = 16'h45b;
#10;
address_ina = 98;
address_inb = 99;
data_ina = 16'h3e0;
data_inb = 16'h128;
#10;
address_ina = 100;
address_inb = 101;
data_ina = 16'h18d;
data_inb = 16'h7b5;
#10;
address_ina = 102;
address_inb = 103;
data_ina = 16'h1d1;
data_inb = 16'h236;
#10;
address_ina = 104;
address_inb = 105;
data_ina = 16'h1a7;
data_inb = 16'h256;
#10;
address_ina = 106;
address_inb = 107;
data_ina = 16'h532;
data_inb = 16'h9c;
#10;
address_ina = 108;
address_inb = 109;
data_ina = 16'h36b;
data_inb = 16'h7c2;
#10;
address_ina = 110;
address_inb = 111;
data_ina = 16'ha40;
data_inb = 16'h781;
#10;
address_ina = 112;
address_inb = 113;
data_ina = 16'h155;
data_inb = 16'h6f;
#10;
address_ina = 114;
address_inb = 115;
data_ina = 16'hc14;
data_inb = 16'ha02;
#10;
address_ina = 116;
address_inb = 117;
data_ina = 16'ha02;
data_inb = 16'haa8;
#10;
address_ina = 118;
address_inb = 119;
data_ina = 16'h24;
data_inb = 16'h53b;
#10;
address_ina = 120;
address_inb = 121;
data_ina = 16'h3;
data_inb = 16'h448;
#10;
address_ina = 122;
address_inb = 123;
data_ina = 16'hc96;
data_inb = 16'h9f5;
#10;
address_ina = 124;
address_inb = 125;
data_ina = 16'h1a3;
data_inb = 16'h6b;
#10;
address_ina = 126;
address_inb = 127;
data_ina = 16'h4f7;
data_inb = 16'h7a8;
#10;
address_ina = 128;
address_inb = 129;
data_ina = 16'hb0;
data_inb = 16'h462;
#10;
address_ina = 130;
address_inb = 131;
data_ina = 16'h229;
data_inb = 16'h781;
#10;
address_ina = 132;
address_inb = 133;
data_ina = 16'h6a4;
data_inb = 16'h8ea;
#10;
address_ina = 134;
address_inb = 135;
data_ina = 16'h761;
data_inb = 16'h851;
#10;
address_ina = 136;
address_inb = 137;
data_ina = 16'hcca;
data_inb = 16'h639;
#10;
address_ina = 138;
address_inb = 139;
data_ina = 16'h34d;
data_inb = 16'h636;
#10;
address_ina = 140;
address_inb = 141;
data_ina = 16'h81a;
data_inb = 16'haa4;
#10;
address_ina = 142;
address_inb = 143;
data_ina = 16'hbdc;
data_inb = 16'h8da;
#10;
address_ina = 144;
address_inb = 145;
data_ina = 16'h514;
data_inb = 16'h848;
#10;
address_ina = 146;
address_inb = 147;
data_ina = 16'ha5d;
data_inb = 16'h9a3;
#10;
address_ina = 148;
address_inb = 149;
data_ina = 16'h421;
data_inb = 16'h969;
#10;
address_ina = 150;
address_inb = 151;
data_ina = 16'hc24;
data_inb = 16'h552;
#10;
address_ina = 152;
address_inb = 153;
data_ina = 16'h925;
data_inb = 16'h36e;
#10;
address_ina = 154;
address_inb = 155;
data_ina = 16'h706;
data_inb = 16'h8a3;
#10;
address_ina = 156;
address_inb = 157;
data_ina = 16'hc3b;
data_inb = 16'h72a;
#10;
address_ina = 158;
address_inb = 159;
data_ina = 16'h16f;
data_inb = 16'h6cf;
#10;
address_ina = 160;
address_inb = 161;
data_ina = 16'h309;
data_inb = 16'h2c1;
#10;
address_ina = 162;
address_inb = 163;
data_ina = 16'h4fa;
data_inb = 16'h1ee;
#10;
address_ina = 164;
address_inb = 165;
data_ina = 16'hd7;
data_inb = 16'h5e4;
#10;
address_ina = 166;
address_inb = 167;
data_ina = 16'hbbf;
data_inb = 16'hac2;
#10;
address_ina = 168;
address_inb = 169;
data_ina = 16'h800;
data_inb = 16'h306;
#10;
address_ina = 170;
address_inb = 171;
data_ina = 16'h1ca;
data_inb = 16'hb92;
#10;
address_ina = 172;
address_inb = 173;
data_ina = 16'h266;
data_inb = 16'h33d;
#10;
address_ina = 174;
address_inb = 175;
data_ina = 16'h78b;
data_inb = 16'h7e9;
#10;
address_ina = 176;
address_inb = 177;
data_ina = 16'h489;
data_inb = 16'h764;
#10;
address_ina = 178;
address_inb = 179;
data_ina = 16'h22c;
data_inb = 16'h576;
#10;
address_ina = 180;
address_inb = 181;
data_ina = 16'hc6f;
data_inb = 16'h1fe;
#10;
address_ina = 182;
address_inb = 183;
data_ina = 16'haa8;
data_inb = 16'h27d;
#10;
address_ina = 184;
address_inb = 185;
data_ina = 16'h583;
data_inb = 16'h9a0;
#10;
address_ina = 186;
address_inb = 187;
data_ina = 16'h1f8;
data_inb = 16'h9cb;
#10;
address_ina = 188;
address_inb = 189;
data_ina = 16'h855;
data_inb = 16'h27;
#10;
address_ina = 190;
address_inb = 191;
data_ina = 16'h7f;
data_inb = 16'h10e;
#10;
address_ina = 192;
address_inb = 193;
data_ina = 16'h61c;
data_inb = 16'h781;
#10;
address_ina = 194;
address_inb = 195;
data_ina = 16'h872;
data_inb = 16'h496;
#10;
address_ina = 196;
address_inb = 197;
data_ina = 16'h2b4;
data_inb = 16'h166;
#10;
address_ina = 198;
address_inb = 199;
data_ina = 16'h1a7;
data_inb = 16'h5a3;
#10;
address_ina = 200;
address_inb = 201;
data_ina = 16'h4b3;
data_inb = 16'h9d8;
#10;
address_ina = 202;
address_inb = 203;
data_ina = 16'h521;
data_inb = 16'h1c4;
#10;
address_ina = 204;
address_inb = 205;
data_ina = 16'h831;
data_inb = 16'ha60;
#10;
address_ina = 206;
address_inb = 207;
data_ina = 16'h46b;
data_inb = 16'h180;
#10;
address_ina = 208;
address_inb = 209;
data_ina = 16'hc07;
data_inb = 16'h986;
#10;
address_ina = 210;
address_inb = 211;
data_ina = 16'hb57;
data_inb = 16'h552;
#10;
address_ina = 212;
address_inb = 213;
data_ina = 16'ha84;
data_inb = 16'h8c;
#10;
address_ina = 214;
address_inb = 215;
data_ina = 16'h78e;
data_inb = 16'h1f1;
#10;
address_ina = 216;
address_inb = 217;
data_ina = 16'h448;
data_inb = 16'h395;
#10;
address_ina = 218;
address_inb = 219;
data_ina = 16'h43e;
data_inb = 16'h528;
#10;
address_ina = 220;
address_inb = 221;
data_ina = 16'h3b2;
data_inb = 16'h183;
#10;
address_ina = 222;
address_inb = 223;
data_ina = 16'hc58;
data_inb = 16'h34d;
#10;
address_ina = 224;
address_inb = 225;
data_ina = 16'h8b9;
data_inb = 16'h76b;
#10;
address_ina = 226;
address_inb = 227;
data_ina = 16'h395;
data_inb = 16'h589;
#10;
address_ina = 228;
address_inb = 229;
data_ina = 16'h180;
data_inb = 16'h2a7;
#10;
address_ina = 230;
address_inb = 231;
data_ina = 16'h6c2;
data_inb = 16'h374;
#10;
address_ina = 232;
address_inb = 233;
data_ina = 16'h76e;
data_inb = 16'h6e9;
#10;
address_ina = 234;
address_inb = 235;
data_ina = 16'h8b9;
data_inb = 16'h3a2;
#10;
address_ina = 236;
address_inb = 237;
data_ina = 16'h176;
data_inb = 16'h88c;
#10;
address_ina = 238;
address_inb = 239;
data_ina = 16'h7f;
data_inb = 16'h670;
#10;
address_ina = 240;
address_inb = 241;
data_ina = 16'hd;
data_inb = 16'h21;
#10;
address_ina = 242;
address_inb = 243;
data_ina = 16'he7;
data_inb = 16'h34d;
#10;
address_ina = 244;
address_inb = 245;
data_ina = 16'h4ca;
data_inb = 16'h7d6;
#10;
address_ina = 246;
address_inb = 247;
data_ina = 16'h507;
data_inb = 16'h834;
#10;
address_ina = 248;
address_inb = 249;
data_ina = 16'hb44;
data_inb = 16'h92b;
#10;
address_ina = 250;
address_inb = 251;
data_ina = 16'h319;
data_inb = 16'h75a;
#10;
address_ina = 252;
address_inb = 253;
data_ina = 16'hba5;
data_inb = 16'h6a1;
#10;
address_ina = 254;
address_inb = 255;
data_ina = 16'h91b;
data_inb = 16'h713;
#10;
        wait(init_done);
        #30
        we = 0;
        // Start processing
         
		  #38000

        start = 0;



//        wait (wr_req);
//		  wait (!wr_req);
//		   rd_req = 1;
		  wait(done);
		  #20000
rd_req = 1;
        #70 
		  start = 1;
		 #80 
wait(rd_empty)
rd_req = 0;

$display("Finished the NTT test Number %d",test_num);
////Begin test number #79//////////////
rst = 1;

//#1000
start = 1;
mode = 1; //NTT 0 // INTT 1

// Reset for a few clock cycles

#1000

rst = 0;
test_num = test_num + 1;
#1000
we = 1;
address_ina = 0;
address_inb = 1;
data_ina = 16'h6f;
data_inb = 16'h22e;
#10;
address_ina = 2;
address_inb = 3;
data_ina = 16'h5b6;
data_inb = 16'h2ff;
#10;
address_ina = 4;
address_inb = 5;
data_ina = 16'hbd;
data_inb = 16'h42c;
#10;
address_ina = 6;
address_inb = 7;
data_ina = 16'hfa09;
data_inb = 16'h13b;
#10;
address_ina = 8;
address_inb = 9;
data_ina = 16'h4cc;
data_inb = 16'hf9a5;
#10;
address_ina = 10;
address_inb = 11;
data_ina = 16'hf9ae;
data_inb = 16'h4ef;
#10;
address_ina = 12;
address_inb = 13;
data_ina = 16'hfdf7;
data_inb = 16'h435;
#10;
address_ina = 14;
address_inb = 15;
data_ina = 16'hf9aa;
data_inb = 16'hff9f;
#10;
address_ina = 16;
address_inb = 17;
data_ina = 16'h4e2;
data_inb = 16'h5a1;
#10;
address_ina = 18;
address_inb = 19;
data_ina = 16'h4a7;
data_inb = 16'h2aa;
#10;
address_ina = 20;
address_inb = 21;
data_ina = 16'h22c;
data_inb = 16'h9e;
#10;
address_ina = 22;
address_inb = 23;
data_ina = 16'h590;
data_inb = 16'h456;
#10;
address_ina = 24;
address_inb = 25;
data_ina = 16'h599;
data_inb = 16'h2d5;
#10;
address_ina = 26;
address_inb = 27;
data_ina = 16'h53b;
data_inb = 16'h420;
#10;
address_ina = 28;
address_inb = 29;
data_ina = 16'h26d;
data_inb = 16'h554;
#10;
address_ina = 30;
address_inb = 31;
data_ina = 16'h122;
data_inb = 16'hff8d;
#10;
address_ina = 32;
address_inb = 33;
data_ina = 16'h40f;
data_inb = 16'hfa40;
#10;
address_ina = 34;
address_inb = 35;
data_ina = 16'hfee9;
data_inb = 16'h24e;
#10;
address_ina = 36;
address_inb = 37;
data_ina = 16'hfe1a;
data_inb = 16'h2eb;
#10;
address_ina = 38;
address_inb = 39;
data_ina = 16'h457;
data_inb = 16'h1f8;
#10;
address_ina = 40;
address_inb = 41;
data_ina = 16'h169;
data_inb = 16'hfe61;
#10;
address_ina = 42;
address_inb = 43;
data_ina = 16'h4c8;
data_inb = 16'hf9ed;
#10;
address_ina = 44;
address_inb = 45;
data_ina = 16'h1fe;
data_inb = 16'hfdaf;
#10;
address_ina = 46;
address_inb = 47;
data_ina = 16'hd6;
data_inb = 16'hfb30;
#10;
address_ina = 48;
address_inb = 49;
data_ina = 16'hfece;
data_inb = 16'hfb22;
#10;
address_ina = 50;
address_inb = 51;
data_ina = 16'hff84;
data_inb = 16'h2a2;
#10;
address_ina = 52;
address_inb = 53;
data_ina = 16'h5e3;
data_inb = 16'hfe7f;
#10;
address_ina = 54;
address_inb = 55;
data_ina = 16'hffbd;
data_inb = 16'h643;
#10;
address_ina = 56;
address_inb = 57;
data_ina = 16'hfdcc;
data_inb = 16'h52a;
#10;
address_ina = 58;
address_inb = 59;
data_ina = 16'hfc9d;
data_inb = 16'hfd2e;
#10;
address_ina = 60;
address_inb = 61;
data_ina = 16'h463;
data_inb = 16'hfcdc;
#10;
address_ina = 62;
address_inb = 63;
data_ina = 16'h3b0;
data_inb = 16'hfe53;
#10;
address_ina = 64;
address_inb = 65;
data_ina = 16'h58b;
data_inb = 16'h63d;
#10;
address_ina = 66;
address_inb = 67;
data_ina = 16'he1;
data_inb = 16'hf98e;
#10;
address_ina = 68;
address_inb = 69;
data_ina = 16'h43c;
data_inb = 16'hfb6c;
#10;
address_ina = 70;
address_inb = 71;
data_ina = 16'hfb4c;
data_inb = 16'h3d4;
#10;
address_ina = 72;
address_inb = 73;
data_ina = 16'hfd7f;
data_inb = 16'h1a;
#10;
address_ina = 74;
address_inb = 75;
data_ina = 16'hfefb;
data_inb = 16'hfe7b;
#10;
address_ina = 76;
address_inb = 77;
data_ina = 16'h4be;
data_inb = 16'h284;
#10;
address_ina = 78;
address_inb = 79;
data_ina = 16'h2f9;
data_inb = 16'hffa6;
#10;
address_ina = 80;
address_inb = 81;
data_ina = 16'hfb5c;
data_inb = 16'h300;
#10;
address_ina = 82;
address_inb = 83;
data_ina = 16'hfdd6;
data_inb = 16'h1b8;
#10;
address_ina = 84;
address_inb = 85;
data_ina = 16'h41b;
data_inb = 16'hfbbc;
#10;
address_ina = 86;
address_inb = 87;
data_ina = 16'hfde1;
data_inb = 16'h389;
#10;
address_ina = 88;
address_inb = 89;
data_ina = 16'h5c3;
data_inb = 16'hfca5;
#10;
address_ina = 90;
address_inb = 91;
data_ina = 16'hfd7c;
data_inb = 16'h76;
#10;
address_ina = 92;
address_inb = 93;
data_ina = 16'h587;
data_inb = 16'hfe9e;
#10;
address_ina = 94;
address_inb = 95;
data_ina = 16'hfd2b;
data_inb = 16'hfed3;
#10;
address_ina = 96;
address_inb = 97;
data_ina = 16'hff1f;
data_inb = 16'h4f6;
#10;
address_ina = 98;
address_inb = 99;
data_ina = 16'hfc34;
data_inb = 16'h1da;
#10;
address_ina = 100;
address_inb = 101;
data_ina = 16'h643;
data_inb = 16'hfb04;
#10;
address_ina = 102;
address_inb = 103;
data_ina = 16'h94;
data_inb = 16'h20b;
#10;
address_ina = 104;
address_inb = 105;
data_ina = 16'h441;
data_inb = 16'hfc02;
#10;
address_ina = 106;
address_inb = 107;
data_ina = 16'h4e6;
data_inb = 16'h5e4;
#10;
address_ina = 108;
address_inb = 109;
data_ina = 16'hfc4f;
data_inb = 16'hf982;
#10;
address_ina = 110;
address_inb = 111;
data_ina = 16'h4bc;
data_inb = 16'hffdb;
#10;
address_ina = 112;
address_inb = 113;
data_ina = 16'hf3;
data_inb = 16'h2e0;
#10;
address_ina = 114;
address_inb = 115;
data_ina = 16'hfea0;
data_inb = 16'hfb95;
#10;
address_ina = 116;
address_inb = 117;
data_ina = 16'hfbc0;
data_inb = 16'h5d6;
#10;
address_ina = 118;
address_inb = 119;
data_ina = 16'hfa7c;
data_inb = 16'h53e;
#10;
address_ina = 120;
address_inb = 121;
data_ina = 16'h3eb;
data_inb = 16'h1b2;
#10;
address_ina = 122;
address_inb = 123;
data_ina = 16'h2bb;
data_inb = 16'hfce9;
#10;
address_ina = 124;
address_inb = 125;
data_ina = 16'hfae8;
data_inb = 16'hfcb2;
#10;
address_ina = 126;
address_inb = 127;
data_ina = 16'hffbf;
data_inb = 16'hf9f6;
#10;
address_ina = 128;
address_inb = 129;
data_ina = 16'h60e;
data_inb = 16'h77;
#10;
address_ina = 130;
address_inb = 131;
data_ina = 16'h568;
data_inb = 16'hfde5;
#10;
address_ina = 132;
address_inb = 133;
data_ina = 16'h3cc;
data_inb = 16'h3bb;
#10;
address_ina = 134;
address_inb = 135;
data_ina = 16'h247;
data_inb = 16'h63b;
#10;
address_ina = 136;
address_inb = 137;
data_ina = 16'hfa08;
data_inb = 16'hfa27;
#10;
address_ina = 138;
address_inb = 139;
data_ina = 16'hfa12;
data_inb = 16'hfe0d;
#10;
address_ina = 140;
address_inb = 141;
data_ina = 16'h5db;
data_inb = 16'h612;
#10;
address_ina = 142;
address_inb = 143;
data_ina = 16'hfa87;
data_inb = 16'h72;
#10;
address_ina = 144;
address_inb = 145;
data_ina = 16'hff1a;
data_inb = 16'h1bd;
#10;
address_ina = 146;
address_inb = 147;
data_ina = 16'h2f0;
data_inb = 16'hfbaa;
#10;
address_ina = 148;
address_inb = 149;
data_ina = 16'h131;
data_inb = 16'h45d;
#10;
address_ina = 150;
address_inb = 151;
data_ina = 16'h62;
data_inb = 16'hfda5;
#10;
address_ina = 152;
address_inb = 153;
data_ina = 16'h14;
data_inb = 16'hfa00;
#10;
address_ina = 154;
address_inb = 155;
data_ina = 16'hff4d;
data_inb = 16'h618;
#10;
address_ina = 156;
address_inb = 157;
data_ina = 16'hffa2;
data_inb = 16'hfead;
#10;
address_ina = 158;
address_inb = 159;
data_ina = 16'hfa33;
data_inb = 16'hfc8b;
#10;
address_ina = 160;
address_inb = 161;
data_ina = 16'h352;
data_inb = 16'h11e;
#10;
address_ina = 162;
address_inb = 163;
data_ina = 16'hfdc6;
data_inb = 16'hfe00;
#10;
address_ina = 164;
address_inb = 165;
data_ina = 16'h210;
data_inb = 16'h2a5;
#10;
address_ina = 166;
address_inb = 167;
data_ina = 16'h57b;
data_inb = 16'hfabd;
#10;
address_ina = 168;
address_inb = 169;
data_ina = 16'h532;
data_inb = 16'hfb38;
#10;
address_ina = 170;
address_inb = 171;
data_ina = 16'h51c;
data_inb = 16'h361;
#10;
address_ina = 172;
address_inb = 173;
data_ina = 16'h406;
data_inb = 16'h50e;
#10;
address_ina = 174;
address_inb = 175;
data_ina = 16'h11b;
data_inb = 16'hfa69;
#10;
address_ina = 176;
address_inb = 177;
data_ina = 16'h374;
data_inb = 16'h57e;
#10;
address_ina = 178;
address_inb = 179;
data_ina = 16'hfd2e;
data_inb = 16'hfe52;
#10;
address_ina = 180;
address_inb = 181;
data_ina = 16'hfaa8;
data_inb = 16'h48;
#10;
address_ina = 182;
address_inb = 183;
data_ina = 16'hfa7d;
data_inb = 16'h26e;
#10;
address_ina = 184;
address_inb = 185;
data_ina = 16'h60f;
data_inb = 16'hffa9;
#10;
address_ina = 186;
address_inb = 187;
data_ina = 16'hffcd;
data_inb = 16'h13d;
#10;
address_ina = 188;
address_inb = 189;
data_ina = 16'h267;
data_inb = 16'h318;
#10;
address_ina = 190;
address_inb = 191;
data_ina = 16'hff94;
data_inb = 16'hfa25;
#10;
address_ina = 192;
address_inb = 193;
data_ina = 16'he2;
data_inb = 16'hfdb8;
#10;
address_ina = 194;
address_inb = 195;
data_ina = 16'hf99e;
data_inb = 16'hfda6;
#10;
address_ina = 196;
address_inb = 197;
data_ina = 16'hfcce;
data_inb = 16'h101;
#10;
address_ina = 198;
address_inb = 199;
data_ina = 16'h105;
data_inb = 16'h2fc;
#10;
address_ina = 200;
address_inb = 201;
data_ina = 16'hfdf2;
data_inb = 16'hfa86;
#10;
address_ina = 202;
address_inb = 203;
data_ina = 16'h22f;
data_inb = 16'hfc6d;
#10;
address_ina = 204;
address_inb = 205;
data_ina = 16'hfcca;
data_inb = 16'hfaf2;
#10;
address_ina = 206;
address_inb = 207;
data_ina = 16'h2a8;
data_inb = 16'h455;
#10;
address_ina = 208;
address_inb = 209;
data_ina = 16'h578;
data_inb = 16'h635;
#10;
address_ina = 210;
address_inb = 211;
data_ina = 16'hfada;
data_inb = 16'hff8b;
#10;
address_ina = 212;
address_inb = 213;
data_ina = 16'hfb4d;
data_inb = 16'hfef5;
#10;
address_ina = 214;
address_inb = 215;
data_ina = 16'hed;
data_inb = 16'h7a;
#10;
address_ina = 216;
address_inb = 217;
data_ina = 16'hfe39;
data_inb = 16'h599;
#10;
address_ina = 218;
address_inb = 219;
data_ina = 16'hfa8b;
data_inb = 16'hf99a;
#10;
address_ina = 220;
address_inb = 221;
data_ina = 16'hfef8;
data_inb = 16'h2d2;
#10;
address_ina = 222;
address_inb = 223;
data_ina = 16'h22d;
data_inb = 16'h29c;
#10;
address_ina = 224;
address_inb = 225;
data_ina = 16'h315;
data_inb = 16'h439;
#10;
address_ina = 226;
address_inb = 227;
data_ina = 16'h633;
data_inb = 16'h446;
#10;
address_ina = 228;
address_inb = 229;
data_ina = 16'hf992;
data_inb = 16'hff39;
#10;
address_ina = 230;
address_inb = 231;
data_ina = 16'h440;
data_inb = 16'hb3;
#10;
address_ina = 232;
address_inb = 233;
data_ina = 16'h266;
data_inb = 16'h53f;
#10;
address_ina = 234;
address_inb = 235;
data_ina = 16'hfa90;
data_inb = 16'hf9a2;
#10;
address_ina = 236;
address_inb = 237;
data_ina = 16'h384;
data_inb = 16'h638;
#10;
address_ina = 238;
address_inb = 239;
data_ina = 16'hfb9b;
data_inb = 16'hfcd2;
#10;
address_ina = 240;
address_inb = 241;
data_ina = 16'hc8;
data_inb = 16'hfcec;
#10;
address_ina = 242;
address_inb = 243;
data_ina = 16'h653;
data_inb = 16'hff67;
#10;
address_ina = 244;
address_inb = 245;
data_ina = 16'h5d;
data_inb = 16'hffdf;
#10;
address_ina = 246;
address_inb = 247;
data_ina = 16'h2d1;
data_inb = 16'hfaa9;
#10;
address_ina = 248;
address_inb = 249;
data_ina = 16'hfb4a;
data_inb = 16'h4de;
#10;
address_ina = 250;
address_inb = 251;
data_ina = 16'hfba6;
data_inb = 16'h29c;
#10;
address_ina = 252;
address_inb = 253;
data_ina = 16'hfd55;
data_inb = 16'h27f;
#10;
address_ina = 254;
address_inb = 255;
data_ina = 16'h5f4;
data_inb = 16'h3df;
#10;
        wait(init_done);
        #30
        we = 0;
        // Start processing
         
		  #38000

        start = 0;



//        wait (wr_req);
//		  wait (!wr_req);
//		   rd_req = 1;
		  wait(done);
		  #20000
rd_req = 1;
        #70 
		  start = 1;
		 #80 
wait(rd_empty)
rd_req = 0;

$display("Finished the NTT test Number %d",test_num);
////Begin test number #80//////////////
rst = 1;

//#1000
start = 1;
mode = 0; //NTT 0 // INTT 1

// Reset for a few clock cycles

#1000

rst = 0;
test_num = test_num + 1;
#1000
we = 1;
address_ina = 0;
address_inb = 1;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 2;
address_inb = 3;
data_ina = 16'h2;
data_inb = 16'hffff;
#10;
address_ina = 4;
address_inb = 5;
data_ina = 16'h2;
data_inb = 16'h2;
#10;
address_ina = 6;
address_inb = 7;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 8;
address_inb = 9;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 10;
address_inb = 11;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 12;
address_inb = 13;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 14;
address_inb = 15;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 16;
address_inb = 17;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 18;
address_inb = 19;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 20;
address_inb = 21;
data_ina = 16'h2;
data_inb = 16'h3;
#10;
address_ina = 22;
address_inb = 23;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 24;
address_inb = 25;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 26;
address_inb = 27;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 28;
address_inb = 29;
data_ina = 16'h2;
data_inb = 16'h1;
#10;
address_ina = 30;
address_inb = 31;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 32;
address_inb = 33;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 34;
address_inb = 35;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 36;
address_inb = 37;
data_ina = 16'hfffd;
data_inb = 16'hfffe;
#10;
address_ina = 38;
address_inb = 39;
data_ina = 16'h2;
data_inb = 16'hffff;
#10;
address_ina = 40;
address_inb = 41;
data_ina = 16'h2;
data_inb = 16'hfffe;
#10;
address_ina = 42;
address_inb = 43;
data_ina = 16'h0;
data_inb = 16'h2;
#10;
address_ina = 44;
address_inb = 45;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 46;
address_inb = 47;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 48;
address_inb = 49;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 50;
address_inb = 51;
data_ina = 16'hfffe;
data_inb = 16'h0;
#10;
address_ina = 52;
address_inb = 53;
data_ina = 16'hffff;
data_inb = 16'hfffd;
#10;
address_ina = 54;
address_inb = 55;
data_ina = 16'h3;
data_inb = 16'h0;
#10;
address_ina = 56;
address_inb = 57;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 58;
address_inb = 59;
data_ina = 16'h1;
data_inb = 16'hfffe;
#10;
address_ina = 60;
address_inb = 61;
data_ina = 16'hfffe;
data_inb = 16'h2;
#10;
address_ina = 62;
address_inb = 63;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 64;
address_inb = 65;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 66;
address_inb = 67;
data_ina = 16'hfffe;
data_inb = 16'h2;
#10;
address_ina = 68;
address_inb = 69;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 70;
address_inb = 71;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 72;
address_inb = 73;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 74;
address_inb = 75;
data_ina = 16'h2;
data_inb = 16'h1;
#10;
address_ina = 76;
address_inb = 77;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 78;
address_inb = 79;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 80;
address_inb = 81;
data_ina = 16'h2;
data_inb = 16'hfffd;
#10;
address_ina = 82;
address_inb = 83;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 84;
address_inb = 85;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 86;
address_inb = 87;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 88;
address_inb = 89;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 90;
address_inb = 91;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 92;
address_inb = 93;
data_ina = 16'h2;
data_inb = 16'h0;
#10;
address_ina = 94;
address_inb = 95;
data_ina = 16'h0;
data_inb = 16'h2;
#10;
address_ina = 96;
address_inb = 97;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 98;
address_inb = 99;
data_ina = 16'h0;
data_inb = 16'hfffe;
#10;
address_ina = 100;
address_inb = 101;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 102;
address_inb = 103;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 104;
address_inb = 105;
data_ina = 16'hffff;
data_inb = 16'h2;
#10;
address_ina = 106;
address_inb = 107;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 108;
address_inb = 109;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 110;
address_inb = 111;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 112;
address_inb = 113;
data_ina = 16'hfffe;
data_inb = 16'h3;
#10;
address_ina = 114;
address_inb = 115;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 116;
address_inb = 117;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 118;
address_inb = 119;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 120;
address_inb = 121;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 122;
address_inb = 123;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 124;
address_inb = 125;
data_ina = 16'h2;
data_inb = 16'hffff;
#10;
address_ina = 126;
address_inb = 127;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 128;
address_inb = 129;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 130;
address_inb = 131;
data_ina = 16'hfffe;
data_inb = 16'hfffd;
#10;
address_ina = 132;
address_inb = 133;
data_ina = 16'h1;
data_inb = 16'h2;
#10;
address_ina = 134;
address_inb = 135;
data_ina = 16'hfffe;
data_inb = 16'hffff;
#10;
address_ina = 136;
address_inb = 137;
data_ina = 16'h3;
data_inb = 16'h2;
#10;
address_ina = 138;
address_inb = 139;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 140;
address_inb = 141;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 142;
address_inb = 143;
data_ina = 16'hffff;
data_inb = 16'h2;
#10;
address_ina = 144;
address_inb = 145;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 146;
address_inb = 147;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 148;
address_inb = 149;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 150;
address_inb = 151;
data_ina = 16'h3;
data_inb = 16'hfffe;
#10;
address_ina = 152;
address_inb = 153;
data_ina = 16'hfffe;
data_inb = 16'h2;
#10;
address_ina = 154;
address_inb = 155;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 156;
address_inb = 157;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 158;
address_inb = 159;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 160;
address_inb = 161;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 162;
address_inb = 163;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 164;
address_inb = 165;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 166;
address_inb = 167;
data_ina = 16'h1;
data_inb = 16'h3;
#10;
address_ina = 168;
address_inb = 169;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 170;
address_inb = 171;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 172;
address_inb = 173;
data_ina = 16'h2;
data_inb = 16'h1;
#10;
address_ina = 174;
address_inb = 175;
data_ina = 16'hfffe;
data_inb = 16'hffff;
#10;
address_ina = 176;
address_inb = 177;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 178;
address_inb = 179;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 180;
address_inb = 181;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 182;
address_inb = 183;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 184;
address_inb = 185;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 186;
address_inb = 187;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 188;
address_inb = 189;
data_ina = 16'hffff;
data_inb = 16'hfffe;
#10;
address_ina = 190;
address_inb = 191;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 192;
address_inb = 193;
data_ina = 16'h2;
data_inb = 16'hffff;
#10;
address_ina = 194;
address_inb = 195;
data_ina = 16'hfffe;
data_inb = 16'h0;
#10;
address_ina = 196;
address_inb = 197;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 198;
address_inb = 199;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 200;
address_inb = 201;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 202;
address_inb = 203;
data_ina = 16'h0;
data_inb = 16'h2;
#10;
address_ina = 204;
address_inb = 205;
data_ina = 16'hfffe;
data_inb = 16'hffff;
#10;
address_ina = 206;
address_inb = 207;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 208;
address_inb = 209;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 210;
address_inb = 211;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 212;
address_inb = 213;
data_ina = 16'h1;
data_inb = 16'hfffd;
#10;
address_ina = 214;
address_inb = 215;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 216;
address_inb = 217;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 218;
address_inb = 219;
data_ina = 16'h0;
data_inb = 16'hfffd;
#10;
address_ina = 220;
address_inb = 221;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 222;
address_inb = 223;
data_ina = 16'hfffd;
data_inb = 16'hffff;
#10;
address_ina = 224;
address_inb = 225;
data_ina = 16'h2;
data_inb = 16'hffff;
#10;
address_ina = 226;
address_inb = 227;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 228;
address_inb = 229;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 230;
address_inb = 231;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 232;
address_inb = 233;
data_ina = 16'h2;
data_inb = 16'h1;
#10;
address_ina = 234;
address_inb = 235;
data_ina = 16'hfffe;
data_inb = 16'h0;
#10;
address_ina = 236;
address_inb = 237;
data_ina = 16'h2;
data_inb = 16'h1;
#10;
address_ina = 238;
address_inb = 239;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 240;
address_inb = 241;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 242;
address_inb = 243;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 244;
address_inb = 245;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 246;
address_inb = 247;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 248;
address_inb = 249;
data_ina = 16'h2;
data_inb = 16'h1;
#10;
address_ina = 250;
address_inb = 251;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 252;
address_inb = 253;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 254;
address_inb = 255;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
        wait(init_done);
        #30
        we = 0;
        // Start processing
         
		  #38000

        start = 0;



//        wait (wr_req);
//		  wait (!wr_req);
//		   rd_req = 1;
		  wait(done);
		  #20000
rd_req = 1;
        #70 
		  start = 1;
		 #80 
wait(rd_empty)
rd_req = 0;

$display("Finished the NTT test Number %d",test_num);
////Begin test number #81//////////////
rst = 1;

//#1000
start = 1;
mode = 0; //NTT 0 // INTT 1

// Reset for a few clock cycles

#1000

rst = 0;
test_num = test_num + 1;
#1000
we = 1;
address_ina = 0;
address_inb = 1;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 2;
address_inb = 3;
data_ina = 16'hfffd;
data_inb = 16'h1;
#10;
address_ina = 4;
address_inb = 5;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 6;
address_inb = 7;
data_ina = 16'hffff;
data_inb = 16'h2;
#10;
address_ina = 8;
address_inb = 9;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 10;
address_inb = 11;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 12;
address_inb = 13;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 14;
address_inb = 15;
data_ina = 16'hfffe;
data_inb = 16'h2;
#10;
address_ina = 16;
address_inb = 17;
data_ina = 16'hffff;
data_inb = 16'hfffe;
#10;
address_ina = 18;
address_inb = 19;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 20;
address_inb = 21;
data_ina = 16'h0;
data_inb = 16'h2;
#10;
address_ina = 22;
address_inb = 23;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 24;
address_inb = 25;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 26;
address_inb = 27;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 28;
address_inb = 29;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 30;
address_inb = 31;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 32;
address_inb = 33;
data_ina = 16'h1;
data_inb = 16'hfffe;
#10;
address_ina = 34;
address_inb = 35;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 36;
address_inb = 37;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 38;
address_inb = 39;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 40;
address_inb = 41;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 42;
address_inb = 43;
data_ina = 16'hffff;
data_inb = 16'h2;
#10;
address_ina = 44;
address_inb = 45;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 46;
address_inb = 47;
data_ina = 16'h0;
data_inb = 16'hfffe;
#10;
address_ina = 48;
address_inb = 49;
data_ina = 16'h0;
data_inb = 16'hfffd;
#10;
address_ina = 50;
address_inb = 51;
data_ina = 16'h0;
data_inb = 16'h2;
#10;
address_ina = 52;
address_inb = 53;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 54;
address_inb = 55;
data_ina = 16'h0;
data_inb = 16'h2;
#10;
address_ina = 56;
address_inb = 57;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 58;
address_inb = 59;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 60;
address_inb = 61;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 62;
address_inb = 63;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 64;
address_inb = 65;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 66;
address_inb = 67;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 68;
address_inb = 69;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 70;
address_inb = 71;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 72;
address_inb = 73;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 74;
address_inb = 75;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 76;
address_inb = 77;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 78;
address_inb = 79;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 80;
address_inb = 81;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 82;
address_inb = 83;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 84;
address_inb = 85;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 86;
address_inb = 87;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 88;
address_inb = 89;
data_ina = 16'hfffe;
data_inb = 16'h1;
#10;
address_ina = 90;
address_inb = 91;
data_ina = 16'h2;
data_inb = 16'h1;
#10;
address_ina = 92;
address_inb = 93;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 94;
address_inb = 95;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 96;
address_inb = 97;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 98;
address_inb = 99;
data_ina = 16'h1;
data_inb = 16'hfffe;
#10;
address_ina = 100;
address_inb = 101;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 102;
address_inb = 103;
data_ina = 16'h0;
data_inb = 16'h2;
#10;
address_ina = 104;
address_inb = 105;
data_ina = 16'hfffe;
data_inb = 16'h1;
#10;
address_ina = 106;
address_inb = 107;
data_ina = 16'h2;
data_inb = 16'hffff;
#10;
address_ina = 108;
address_inb = 109;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 110;
address_inb = 111;
data_ina = 16'h3;
data_inb = 16'h0;
#10;
address_ina = 112;
address_inb = 113;
data_ina = 16'h1;
data_inb = 16'h2;
#10;
address_ina = 114;
address_inb = 115;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 116;
address_inb = 117;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 118;
address_inb = 119;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 120;
address_inb = 121;
data_ina = 16'h3;
data_inb = 16'hfffe;
#10;
address_ina = 122;
address_inb = 123;
data_ina = 16'h0;
data_inb = 16'h2;
#10;
address_ina = 124;
address_inb = 125;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 126;
address_inb = 127;
data_ina = 16'h2;
data_inb = 16'hffff;
#10;
address_ina = 128;
address_inb = 129;
data_ina = 16'h2;
data_inb = 16'hffff;
#10;
address_ina = 130;
address_inb = 131;
data_ina = 16'h2;
data_inb = 16'hfffd;
#10;
address_ina = 132;
address_inb = 133;
data_ina = 16'h3;
data_inb = 16'h0;
#10;
address_ina = 134;
address_inb = 135;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 136;
address_inb = 137;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 138;
address_inb = 139;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 140;
address_inb = 141;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 142;
address_inb = 143;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 144;
address_inb = 145;
data_ina = 16'h1;
data_inb = 16'h2;
#10;
address_ina = 146;
address_inb = 147;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 148;
address_inb = 149;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 150;
address_inb = 151;
data_ina = 16'hfffe;
data_inb = 16'hffff;
#10;
address_ina = 152;
address_inb = 153;
data_ina = 16'hfffe;
data_inb = 16'h2;
#10;
address_ina = 154;
address_inb = 155;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 156;
address_inb = 157;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 158;
address_inb = 159;
data_ina = 16'hfffe;
data_inb = 16'h1;
#10;
address_ina = 160;
address_inb = 161;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 162;
address_inb = 163;
data_ina = 16'hfffe;
data_inb = 16'hfffe;
#10;
address_ina = 164;
address_inb = 165;
data_ina = 16'h2;
data_inb = 16'h2;
#10;
address_ina = 166;
address_inb = 167;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 168;
address_inb = 169;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 170;
address_inb = 171;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 172;
address_inb = 173;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 174;
address_inb = 175;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 176;
address_inb = 177;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 178;
address_inb = 179;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 180;
address_inb = 181;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 182;
address_inb = 183;
data_ina = 16'h0;
data_inb = 16'hfffe;
#10;
address_ina = 184;
address_inb = 185;
data_ina = 16'h0;
data_inb = 16'h2;
#10;
address_ina = 186;
address_inb = 187;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 188;
address_inb = 189;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 190;
address_inb = 191;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 192;
address_inb = 193;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 194;
address_inb = 195;
data_ina = 16'h2;
data_inb = 16'h1;
#10;
address_ina = 196;
address_inb = 197;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 198;
address_inb = 199;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 200;
address_inb = 201;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 202;
address_inb = 203;
data_ina = 16'hfffd;
data_inb = 16'h1;
#10;
address_ina = 204;
address_inb = 205;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 206;
address_inb = 207;
data_ina = 16'h0;
data_inb = 16'hfffe;
#10;
address_ina = 208;
address_inb = 209;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 210;
address_inb = 211;
data_ina = 16'hfffe;
data_inb = 16'hffff;
#10;
address_ina = 212;
address_inb = 213;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 214;
address_inb = 215;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 216;
address_inb = 217;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 218;
address_inb = 219;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 220;
address_inb = 221;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 222;
address_inb = 223;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 224;
address_inb = 225;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 226;
address_inb = 227;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 228;
address_inb = 229;
data_ina = 16'hfffe;
data_inb = 16'h0;
#10;
address_ina = 230;
address_inb = 231;
data_ina = 16'h0;
data_inb = 16'h2;
#10;
address_ina = 232;
address_inb = 233;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 234;
address_inb = 235;
data_ina = 16'h1;
data_inb = 16'hfffe;
#10;
address_ina = 236;
address_inb = 237;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 238;
address_inb = 239;
data_ina = 16'hfffe;
data_inb = 16'h1;
#10;
address_ina = 240;
address_inb = 241;
data_ina = 16'h0;
data_inb = 16'hfffe;
#10;
address_ina = 242;
address_inb = 243;
data_ina = 16'h3;
data_inb = 16'h0;
#10;
address_ina = 244;
address_inb = 245;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 246;
address_inb = 247;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 248;
address_inb = 249;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 250;
address_inb = 251;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 252;
address_inb = 253;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 254;
address_inb = 255;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
        wait(init_done);
        #30
        we = 0;
        // Start processing
         
		  #38000

        start = 0;



//        wait (wr_req);
//		  wait (!wr_req);
//		   rd_req = 1;
		  wait(done);
		  #20000
rd_req = 1;
        #70 
		  start = 1;
		 #80 
wait(rd_empty)
rd_req = 0;

$display("Finished the NTT test Number %d",test_num);
////Begin test number #82//////////////
rst = 1;

//#1000
start = 1;
mode = 1; //NTT 0 // INTT 1

// Reset for a few clock cycles

#1000

rst = 0;
test_num = test_num + 1;
#1000
we = 1;
address_ina = 0;
address_inb = 1;
data_ina = 16'hfc39;
data_inb = 16'hff11;
#10;
address_ina = 2;
address_inb = 3;
data_ina = 16'hfd0a;
data_inb = 16'hfcda;
#10;
address_ina = 4;
address_inb = 5;
data_ina = 16'h2fa;
data_inb = 16'hfdbf;
#10;
address_ina = 6;
address_inb = 7;
data_ina = 16'h5f6;
data_inb = 16'hfc5c;
#10;
address_ina = 8;
address_inb = 9;
data_ina = 16'h1e5;
data_inb = 16'hfbe9;
#10;
address_ina = 10;
address_inb = 11;
data_ina = 16'h45e;
data_inb = 16'hfc6b;
#10;
address_ina = 12;
address_inb = 13;
data_ina = 16'h573;
data_inb = 16'h515;
#10;
address_ina = 14;
address_inb = 15;
data_ina = 16'hfa39;
data_inb = 16'hf9d6;
#10;
address_ina = 16;
address_inb = 17;
data_ina = 16'h2d7;
data_inb = 16'hfd8f;
#10;
address_ina = 18;
address_inb = 19;
data_ina = 16'h401;
data_inb = 16'hfa45;
#10;
address_ina = 20;
address_inb = 21;
data_ina = 16'hfbd1;
data_inb = 16'hfa78;
#10;
address_ina = 22;
address_inb = 23;
data_ina = 16'hff14;
data_inb = 16'h1c7;
#10;
address_ina = 24;
address_inb = 25;
data_ina = 16'h4a7;
data_inb = 16'hfdd5;
#10;
address_ina = 26;
address_inb = 27;
data_ina = 16'hf9b4;
data_inb = 16'hff41;
#10;
address_ina = 28;
address_inb = 29;
data_ina = 16'h5e0;
data_inb = 16'hfc42;
#10;
address_ina = 30;
address_inb = 31;
data_ina = 16'hfc55;
data_inb = 16'h399;
#10;
address_ina = 32;
address_inb = 33;
data_ina = 16'h658;
data_inb = 16'h1af;
#10;
address_ina = 34;
address_inb = 35;
data_ina = 16'hfa9e;
data_inb = 16'h1bc;
#10;
address_ina = 36;
address_inb = 37;
data_ina = 16'h4ac;
data_inb = 16'hfbc7;
#10;
address_ina = 38;
address_inb = 39;
data_ina = 16'h5e6;
data_inb = 16'h460;
#10;
address_ina = 40;
address_inb = 41;
data_ina = 16'hfea4;
data_inb = 16'h367;
#10;
address_ina = 42;
address_inb = 43;
data_ina = 16'hfa35;
data_inb = 16'h235;
#10;
address_ina = 44;
address_inb = 45;
data_ina = 16'h43f;
data_inb = 16'h14f;
#10;
address_ina = 46;
address_inb = 47;
data_ina = 16'hfe7c;
data_inb = 16'hfed2;
#10;
address_ina = 48;
address_inb = 49;
data_ina = 16'hff5f;
data_inb = 16'hfe3a;
#10;
address_ina = 50;
address_inb = 51;
data_ina = 16'h524;
data_inb = 16'h81;
#10;
address_ina = 52;
address_inb = 53;
data_ina = 16'h5ef;
data_inb = 16'h2e0;
#10;
address_ina = 54;
address_inb = 55;
data_ina = 16'hfb00;
data_inb = 16'hfa25;
#10;
address_ina = 56;
address_inb = 57;
data_ina = 16'hfc70;
data_inb = 16'hfc16;
#10;
address_ina = 58;
address_inb = 59;
data_ina = 16'h3a1;
data_inb = 16'hfe1d;
#10;
address_ina = 60;
address_inb = 61;
data_ina = 16'hfd07;
data_inb = 16'h8b;
#10;
address_ina = 62;
address_inb = 63;
data_ina = 16'hfed1;
data_inb = 16'h3a;
#10;
address_ina = 64;
address_inb = 65;
data_ina = 16'h1ec;
data_inb = 16'h2f5;
#10;
address_ina = 66;
address_inb = 67;
data_ina = 16'h5f7;
data_inb = 16'hfd20;
#10;
address_ina = 68;
address_inb = 69;
data_ina = 16'h665;
data_inb = 16'h457;
#10;
address_ina = 70;
address_inb = 71;
data_ina = 16'hfba9;
data_inb = 16'hfbc9;
#10;
address_ina = 72;
address_inb = 73;
data_ina = 16'hffd5;
data_inb = 16'hfd73;
#10;
address_ina = 74;
address_inb = 75;
data_ina = 16'h2ef;
data_inb = 16'hfcd7;
#10;
address_ina = 76;
address_inb = 77;
data_ina = 16'hff0d;
data_inb = 16'hfd4c;
#10;
address_ina = 78;
address_inb = 79;
data_ina = 16'h15e;
data_inb = 16'hfdf8;
#10;
address_ina = 80;
address_inb = 81;
data_ina = 16'hfcf4;
data_inb = 16'hfa33;
#10;
address_ina = 82;
address_inb = 83;
data_ina = 16'h4d6;
data_inb = 16'hfa14;
#10;
address_ina = 84;
address_inb = 85;
data_ina = 16'hd3;
data_inb = 16'hfa16;
#10;
address_ina = 86;
address_inb = 87;
data_ina = 16'hfd2f;
data_inb = 16'h24d;
#10;
address_ina = 88;
address_inb = 89;
data_ina = 16'hfe3c;
data_inb = 16'hfcec;
#10;
address_ina = 90;
address_inb = 91;
data_ina = 16'h35e;
data_inb = 16'h10e;
#10;
address_ina = 92;
address_inb = 93;
data_ina = 16'h16a;
data_inb = 16'h2f;
#10;
address_ina = 94;
address_inb = 95;
data_ina = 16'hfc9e;
data_inb = 16'h1b7;
#10;
address_ina = 96;
address_inb = 97;
data_ina = 16'h374;
data_inb = 16'h33f;
#10;
address_ina = 98;
address_inb = 99;
data_ina = 16'h407;
data_inb = 16'hff7d;
#10;
address_ina = 100;
address_inb = 101;
data_ina = 16'hff3f;
data_inb = 16'hfde7;
#10;
address_ina = 102;
address_inb = 103;
data_ina = 16'h4b;
data_inb = 16'h155;
#10;
address_ina = 104;
address_inb = 105;
data_ina = 16'hff6b;
data_inb = 16'hfc;
#10;
address_ina = 106;
address_inb = 107;
data_ina = 16'h375;
data_inb = 16'hfc79;
#10;
address_ina = 108;
address_inb = 109;
data_ina = 16'hfb41;
data_inb = 16'h101;
#10;
address_ina = 110;
address_inb = 111;
data_ina = 16'hfd6c;
data_inb = 16'hfa95;
#10;
address_ina = 112;
address_inb = 113;
data_ina = 16'h664;
data_inb = 16'h395;
#10;
address_ina = 114;
address_inb = 115;
data_ina = 16'h46d;
data_inb = 16'hfe89;
#10;
address_ina = 116;
address_inb = 117;
data_ina = 16'hfce3;
data_inb = 16'hfa4e;
#10;
address_ina = 118;
address_inb = 119;
data_ina = 16'h663;
data_inb = 16'hfd51;
#10;
address_ina = 120;
address_inb = 121;
data_ina = 16'hfe3e;
data_inb = 16'hfdee;
#10;
address_ina = 122;
address_inb = 123;
data_ina = 16'h311;
data_inb = 16'hfe51;
#10;
address_ina = 124;
address_inb = 125;
data_ina = 16'hfdfc;
data_inb = 16'hff35;
#10;
address_ina = 126;
address_inb = 127;
data_ina = 16'h29b;
data_inb = 16'h531;
#10;
address_ina = 128;
address_inb = 129;
data_ina = 16'hfe83;
data_inb = 16'hf9a8;
#10;
address_ina = 130;
address_inb = 131;
data_ina = 16'hffe1;
data_inb = 16'hfb98;
#10;
address_ina = 132;
address_inb = 133;
data_ina = 16'hfd99;
data_inb = 16'h651;
#10;
address_ina = 134;
address_inb = 135;
data_ina = 16'h3fb;
data_inb = 16'h1f4;
#10;
address_ina = 136;
address_inb = 137;
data_ina = 16'h298;
data_inb = 16'hfb10;
#10;
address_ina = 138;
address_inb = 139;
data_ina = 16'hfb4d;
data_inb = 16'hfc42;
#10;
address_ina = 140;
address_inb = 141;
data_ina = 16'hfcf2;
data_inb = 16'hfd51;
#10;
address_ina = 142;
address_inb = 143;
data_ina = 16'hffb1;
data_inb = 16'h61c;
#10;
address_ina = 144;
address_inb = 145;
data_ina = 16'h525;
data_inb = 16'hfa8c;
#10;
address_ina = 146;
address_inb = 147;
data_ina = 16'hfaa9;
data_inb = 16'h1b8;
#10;
address_ina = 148;
address_inb = 149;
data_ina = 16'h323;
data_inb = 16'h43c;
#10;
address_ina = 150;
address_inb = 151;
data_ina = 16'hfa30;
data_inb = 16'he3;
#10;
address_ina = 152;
address_inb = 153;
data_ina = 16'h424;
data_inb = 16'hfeba;
#10;
address_ina = 154;
address_inb = 155;
data_ina = 16'hfbd8;
data_inb = 16'h22f;
#10;
address_ina = 156;
address_inb = 157;
data_ina = 16'hfe3e;
data_inb = 16'hfd53;
#10;
address_ina = 158;
address_inb = 159;
data_ina = 16'hfda5;
data_inb = 16'hfbe1;
#10;
address_ina = 160;
address_inb = 161;
data_ina = 16'hfc77;
data_inb = 16'h5f4;
#10;
address_ina = 162;
address_inb = 163;
data_ina = 16'hfe74;
data_inb = 16'hfbf9;
#10;
address_ina = 164;
address_inb = 165;
data_ina = 16'h3ba;
data_inb = 16'h438;
#10;
address_ina = 166;
address_inb = 167;
data_ina = 16'h5ef;
data_inb = 16'hfdf1;
#10;
address_ina = 168;
address_inb = 169;
data_ina = 16'h1d0;
data_inb = 16'h636;
#10;
address_ina = 170;
address_inb = 171;
data_ina = 16'h119;
data_inb = 16'hfba5;
#10;
address_ina = 172;
address_inb = 173;
data_ina = 16'hfbbc;
data_inb = 16'hffe3;
#10;
address_ina = 174;
address_inb = 175;
data_ina = 16'h486;
data_inb = 16'hfe;
#10;
address_ina = 176;
address_inb = 177;
data_ina = 16'hfd46;
data_inb = 16'hfc45;
#10;
address_ina = 178;
address_inb = 179;
data_ina = 16'h341;
data_inb = 16'hf990;
#10;
address_ina = 180;
address_inb = 181;
data_ina = 16'hab;
data_inb = 16'hf9d6;
#10;
address_ina = 182;
address_inb = 183;
data_ina = 16'hfb4f;
data_inb = 16'hfc95;
#10;
address_ina = 184;
address_inb = 185;
data_ina = 16'h1;
data_inb = 16'hf9b5;
#10;
address_ina = 186;
address_inb = 187;
data_ina = 16'h1e0;
data_inb = 16'hfa64;
#10;
address_ina = 188;
address_inb = 189;
data_ina = 16'h4da;
data_inb = 16'h3b0;
#10;
address_ina = 190;
address_inb = 191;
data_ina = 16'h207;
data_inb = 16'h7b;
#10;
address_ina = 192;
address_inb = 193;
data_ina = 16'h381;
data_inb = 16'hfbcb;
#10;
address_ina = 194;
address_inb = 195;
data_ina = 16'hfd94;
data_inb = 16'hfd17;
#10;
address_ina = 196;
address_inb = 197;
data_ina = 16'h62b;
data_inb = 16'hfd71;
#10;
address_ina = 198;
address_inb = 199;
data_ina = 16'h1a4;
data_inb = 16'h4f5;
#10;
address_ina = 200;
address_inb = 201;
data_ina = 16'hfe5f;
data_inb = 16'hfb82;
#10;
address_ina = 202;
address_inb = 203;
data_ina = 16'hfb89;
data_inb = 16'h3cd;
#10;
address_ina = 204;
address_inb = 205;
data_ina = 16'h46a;
data_inb = 16'h463;
#10;
address_ina = 206;
address_inb = 207;
data_ina = 16'hff4f;
data_inb = 16'h525;
#10;
address_ina = 208;
address_inb = 209;
data_ina = 16'hba;
data_inb = 16'hf9fa;
#10;
address_ina = 210;
address_inb = 211;
data_ina = 16'h172;
data_inb = 16'hd6;
#10;
address_ina = 212;
address_inb = 213;
data_ina = 16'hffcf;
data_inb = 16'hfb1f;
#10;
address_ina = 214;
address_inb = 215;
data_ina = 16'hfcb1;
data_inb = 16'hfce6;
#10;
address_ina = 216;
address_inb = 217;
data_ina = 16'h265;
data_inb = 16'h52c;
#10;
address_ina = 218;
address_inb = 219;
data_ina = 16'hffbc;
data_inb = 16'hf99c;
#10;
address_ina = 220;
address_inb = 221;
data_ina = 16'h60f;
data_inb = 16'hfcb5;
#10;
address_ina = 222;
address_inb = 223;
data_ina = 16'h424;
data_inb = 16'h2ee;
#10;
address_ina = 224;
address_inb = 225;
data_ina = 16'hfe4a;
data_inb = 16'hfeda;
#10;
address_ina = 226;
address_inb = 227;
data_ina = 16'hf9e9;
data_inb = 16'h477;
#10;
address_ina = 228;
address_inb = 229;
data_ina = 16'h120;
data_inb = 16'hfeb5;
#10;
address_ina = 230;
address_inb = 231;
data_ina = 16'hfa3e;
data_inb = 16'hffd5;
#10;
address_ina = 232;
address_inb = 233;
data_ina = 16'hff13;
data_inb = 16'hfdfa;
#10;
address_ina = 234;
address_inb = 235;
data_ina = 16'hfabd;
data_inb = 16'h312;
#10;
address_ina = 236;
address_inb = 237;
data_ina = 16'hfcdc;
data_inb = 16'hff8a;
#10;
address_ina = 238;
address_inb = 239;
data_ina = 16'h2df;
data_inb = 16'hfdc7;
#10;
address_ina = 240;
address_inb = 241;
data_ina = 16'ha;
data_inb = 16'h41f;
#10;
address_ina = 242;
address_inb = 243;
data_ina = 16'h279;
data_inb = 16'h397;
#10;
address_ina = 244;
address_inb = 245;
data_ina = 16'h167;
data_inb = 16'h222;
#10;
address_ina = 246;
address_inb = 247;
data_ina = 16'hf9ea;
data_inb = 16'h330;
#10;
address_ina = 248;
address_inb = 249;
data_ina = 16'hfe67;
data_inb = 16'h57f;
#10;
address_ina = 250;
address_inb = 251;
data_ina = 16'hff14;
data_inb = 16'hbf;
#10;
address_ina = 252;
address_inb = 253;
data_ina = 16'h248;
data_inb = 16'hfb90;
#10;
address_ina = 254;
address_inb = 255;
data_ina = 16'hfdd6;
data_inb = 16'h3d6;
#10;
        wait(init_done);
        #30
        we = 0;
        // Start processing
         
		  #38000

        start = 0;



//        wait (wr_req);
//		  wait (!wr_req);
//		   rd_req = 1;
		  wait(done);
		  #20000
rd_req = 1;
        #70 
		  start = 1;
		 #80 
wait(rd_empty)
rd_req = 0;

$display("Finished the NTT test Number %d",test_num);
////Begin test number #83//////////////
rst = 1;

//#1000
start = 1;
mode = 1; //NTT 0 // INTT 1

// Reset for a few clock cycles

#1000

rst = 0;
test_num = test_num + 1;
#1000
we = 1;
address_ina = 0;
address_inb = 1;
data_ina = 16'hfb68;
data_inb = 16'h475;
#10;
address_ina = 2;
address_inb = 3;
data_ina = 16'hfbd0;
data_inb = 16'hff3a;
#10;
address_ina = 4;
address_inb = 5;
data_ina = 16'h49;
data_inb = 16'h331;
#10;
address_ina = 6;
address_inb = 7;
data_ina = 16'hfd29;
data_inb = 16'hfca6;
#10;
address_ina = 8;
address_inb = 9;
data_ina = 16'h5fd;
data_inb = 16'hfb1a;
#10;
address_ina = 10;
address_inb = 11;
data_ina = 16'h94;
data_inb = 16'hfc1d;
#10;
address_ina = 12;
address_inb = 13;
data_ina = 16'h1e9;
data_inb = 16'h381;
#10;
address_ina = 14;
address_inb = 15;
data_ina = 16'hfd80;
data_inb = 16'h2f5;
#10;
address_ina = 16;
address_inb = 17;
data_ina = 16'hffee;
data_inb = 16'h41d;
#10;
address_ina = 18;
address_inb = 19;
data_ina = 16'hfac4;
data_inb = 16'h5fc;
#10;
address_ina = 20;
address_inb = 21;
data_ina = 16'hfe7a;
data_inb = 16'hf9ac;
#10;
address_ina = 22;
address_inb = 23;
data_ina = 16'hfa22;
data_inb = 16'h3d6;
#10;
address_ina = 24;
address_inb = 25;
data_ina = 16'h316;
data_inb = 16'h4e0;
#10;
address_ina = 26;
address_inb = 27;
data_ina = 16'h15e;
data_inb = 16'hfe1f;
#10;
address_ina = 28;
address_inb = 29;
data_ina = 16'hfb09;
data_inb = 16'hff62;
#10;
address_ina = 30;
address_inb = 31;
data_ina = 16'hfb64;
data_inb = 16'h182;
#10;
address_ina = 32;
address_inb = 33;
data_ina = 16'h43b;
data_inb = 16'hfda9;
#10;
address_ina = 34;
address_inb = 35;
data_ina = 16'h5b;
data_inb = 16'h2e5;
#10;
address_ina = 36;
address_inb = 37;
data_ina = 16'hfc95;
data_inb = 16'hfca1;
#10;
address_ina = 38;
address_inb = 39;
data_ina = 16'hfc32;
data_inb = 16'hfcf9;
#10;
address_ina = 40;
address_inb = 41;
data_ina = 16'hfa17;
data_inb = 16'h32;
#10;
address_ina = 42;
address_inb = 43;
data_ina = 16'h491;
data_inb = 16'hfe84;
#10;
address_ina = 44;
address_inb = 45;
data_ina = 16'hfe5e;
data_inb = 16'hfdc2;
#10;
address_ina = 46;
address_inb = 47;
data_ina = 16'hfac1;
data_inb = 16'hff39;
#10;
address_ina = 48;
address_inb = 49;
data_ina = 16'h452;
data_inb = 16'h27f;
#10;
address_ina = 50;
address_inb = 51;
data_ina = 16'h2be;
data_inb = 16'h369;
#10;
address_ina = 52;
address_inb = 53;
data_ina = 16'h644;
data_inb = 16'h3ed;
#10;
address_ina = 54;
address_inb = 55;
data_ina = 16'h620;
data_inb = 16'h4c6;
#10;
address_ina = 56;
address_inb = 57;
data_ina = 16'h520;
data_inb = 16'hfa27;
#10;
address_ina = 58;
address_inb = 59;
data_ina = 16'hfba7;
data_inb = 16'hfe68;
#10;
address_ina = 60;
address_inb = 61;
data_ina = 16'hfdcc;
data_inb = 16'hffd6;
#10;
address_ina = 62;
address_inb = 63;
data_ina = 16'h13a;
data_inb = 16'hfcd7;
#10;
address_ina = 64;
address_inb = 65;
data_ina = 16'hfe9e;
data_inb = 16'h3c9;
#10;
address_ina = 66;
address_inb = 67;
data_ina = 16'hfcb6;
data_inb = 16'hfc16;
#10;
address_ina = 68;
address_inb = 69;
data_ina = 16'h268;
data_inb = 16'h526;
#10;
address_ina = 70;
address_inb = 71;
data_ina = 16'h5ea;
data_inb = 16'hfc29;
#10;
address_ina = 72;
address_inb = 73;
data_ina = 16'hfb0a;
data_inb = 16'hac;
#10;
address_ina = 74;
address_inb = 75;
data_ina = 16'hfcc7;
data_inb = 16'h88;
#10;
address_ina = 76;
address_inb = 77;
data_ina = 16'hff09;
data_inb = 16'hfbdd;
#10;
address_ina = 78;
address_inb = 79;
data_ina = 16'h556;
data_inb = 16'h417;
#10;
address_ina = 80;
address_inb = 81;
data_ina = 16'hf9a6;
data_inb = 16'hfb9b;
#10;
address_ina = 82;
address_inb = 83;
data_ina = 16'h407;
data_inb = 16'h44e;
#10;
address_ina = 84;
address_inb = 85;
data_ina = 16'h329;
data_inb = 16'h264;
#10;
address_ina = 86;
address_inb = 87;
data_ina = 16'h46e;
data_inb = 16'h4e8;
#10;
address_ina = 88;
address_inb = 89;
data_ina = 16'hfcb8;
data_inb = 16'h678;
#10;
address_ina = 90;
address_inb = 91;
data_ina = 16'hffe7;
data_inb = 16'hfed2;
#10;
address_ina = 92;
address_inb = 93;
data_ina = 16'hfb18;
data_inb = 16'h338;
#10;
address_ina = 94;
address_inb = 95;
data_ina = 16'hfd16;
data_inb = 16'hfd12;
#10;
address_ina = 96;
address_inb = 97;
data_ina = 16'hfb9d;
data_inb = 16'h2f7;
#10;
address_ina = 98;
address_inb = 99;
data_ina = 16'h1d3;
data_inb = 16'h51c;
#10;
address_ina = 100;
address_inb = 101;
data_ina = 16'hfe93;
data_inb = 16'hfb5e;
#10;
address_ina = 102;
address_inb = 103;
data_ina = 16'hfa98;
data_inb = 16'h94;
#10;
address_ina = 104;
address_inb = 105;
data_ina = 16'hfc87;
data_inb = 16'hfa54;
#10;
address_ina = 106;
address_inb = 107;
data_ina = 16'hf9a9;
data_inb = 16'hfd36;
#10;
address_ina = 108;
address_inb = 109;
data_ina = 16'hfc7b;
data_inb = 16'hfb87;
#10;
address_ina = 110;
address_inb = 111;
data_ina = 16'h638;
data_inb = 16'h606;
#10;
address_ina = 112;
address_inb = 113;
data_ina = 16'h11e;
data_inb = 16'h15e;
#10;
address_ina = 114;
address_inb = 115;
data_ina = 16'h3a1;
data_inb = 16'hfdda;
#10;
address_ina = 116;
address_inb = 117;
data_ina = 16'hfd5b;
data_inb = 16'hc0;
#10;
address_ina = 118;
address_inb = 119;
data_ina = 16'h517;
data_inb = 16'hfc79;
#10;
address_ina = 120;
address_inb = 121;
data_ina = 16'h15c;
data_inb = 16'hfe35;
#10;
address_ina = 122;
address_inb = 123;
data_ina = 16'h4af;
data_inb = 16'hfac6;
#10;
address_ina = 124;
address_inb = 125;
data_ina = 16'h412;
data_inb = 16'hff68;
#10;
address_ina = 126;
address_inb = 127;
data_ina = 16'hf9ab;
data_inb = 16'hfc42;
#10;
address_ina = 128;
address_inb = 129;
data_ina = 16'h3c3;
data_inb = 16'hfc0b;
#10;
address_ina = 130;
address_inb = 131;
data_ina = 16'h502;
data_inb = 16'hff66;
#10;
address_ina = 132;
address_inb = 133;
data_ina = 16'hfa02;
data_inb = 16'hfb5e;
#10;
address_ina = 134;
address_inb = 135;
data_ina = 16'hfb0f;
data_inb = 16'h579;
#10;
address_ina = 136;
address_inb = 137;
data_ina = 16'hfc4f;
data_inb = 16'h59e;
#10;
address_ina = 138;
address_inb = 139;
data_ina = 16'h4c7;
data_inb = 16'hfad7;
#10;
address_ina = 140;
address_inb = 141;
data_ina = 16'hfc02;
data_inb = 16'h348;
#10;
address_ina = 142;
address_inb = 143;
data_ina = 16'hfc4b;
data_inb = 16'hfe3d;
#10;
address_ina = 144;
address_inb = 145;
data_ina = 16'h294;
data_inb = 16'hfb02;
#10;
address_ina = 146;
address_inb = 147;
data_ina = 16'hface;
data_inb = 16'hfcaf;
#10;
address_ina = 148;
address_inb = 149;
data_ina = 16'h4aa;
data_inb = 16'h493;
#10;
address_ina = 150;
address_inb = 151;
data_ina = 16'h70;
data_inb = 16'h2ec;
#10;
address_ina = 152;
address_inb = 153;
data_ina = 16'hfce9;
data_inb = 16'hfeb6;
#10;
address_ina = 154;
address_inb = 155;
data_ina = 16'h1cf;
data_inb = 16'hfdf3;
#10;
address_ina = 156;
address_inb = 157;
data_ina = 16'hfc61;
data_inb = 16'h13b;
#10;
address_ina = 158;
address_inb = 159;
data_ina = 16'hfb2f;
data_inb = 16'h368;
#10;
address_ina = 160;
address_inb = 161;
data_ina = 16'h521;
data_inb = 16'h3c6;
#10;
address_ina = 162;
address_inb = 163;
data_ina = 16'h4af;
data_inb = 16'h118;
#10;
address_ina = 164;
address_inb = 165;
data_ina = 16'hfcc0;
data_inb = 16'hfa3d;
#10;
address_ina = 166;
address_inb = 167;
data_ina = 16'hfae6;
data_inb = 16'hbd;
#10;
address_ina = 168;
address_inb = 169;
data_ina = 16'h314;
data_inb = 16'h51f;
#10;
address_ina = 170;
address_inb = 171;
data_ina = 16'hfbce;
data_inb = 16'hfa4b;
#10;
address_ina = 172;
address_inb = 173;
data_ina = 16'hffa4;
data_inb = 16'h19d;
#10;
address_ina = 174;
address_inb = 175;
data_ina = 16'hf9f0;
data_inb = 16'hfec9;
#10;
address_ina = 176;
address_inb = 177;
data_ina = 16'hf9c7;
data_inb = 16'h476;
#10;
address_ina = 178;
address_inb = 179;
data_ina = 16'hfd20;
data_inb = 16'h30f;
#10;
address_ina = 180;
address_inb = 181;
data_ina = 16'hfaa5;
data_inb = 16'hfcf6;
#10;
address_ina = 182;
address_inb = 183;
data_ina = 16'h467;
data_inb = 16'hfeef;
#10;
address_ina = 184;
address_inb = 185;
data_ina = 16'hfbf7;
data_inb = 16'hfe9f;
#10;
address_ina = 186;
address_inb = 187;
data_ina = 16'h333;
data_inb = 16'hf999;
#10;
address_ina = 188;
address_inb = 189;
data_ina = 16'hfe7b;
data_inb = 16'h128;
#10;
address_ina = 190;
address_inb = 191;
data_ina = 16'hfab4;
data_inb = 16'hfd70;
#10;
address_ina = 192;
address_inb = 193;
data_ina = 16'hfb09;
data_inb = 16'h211;
#10;
address_ina = 194;
address_inb = 195;
data_ina = 16'hfc49;
data_inb = 16'h5dc;
#10;
address_ina = 196;
address_inb = 197;
data_ina = 16'hfd47;
data_inb = 16'h39;
#10;
address_ina = 198;
address_inb = 199;
data_ina = 16'h665;
data_inb = 16'h2f2;
#10;
address_ina = 200;
address_inb = 201;
data_ina = 16'hffb7;
data_inb = 16'h452;
#10;
address_ina = 202;
address_inb = 203;
data_ina = 16'h380;
data_inb = 16'hfbaa;
#10;
address_ina = 204;
address_inb = 205;
data_ina = 16'hfb89;
data_inb = 16'h459;
#10;
address_ina = 206;
address_inb = 207;
data_ina = 16'hfe1a;
data_inb = 16'h19f;
#10;
address_ina = 208;
address_inb = 209;
data_ina = 16'h55a;
data_inb = 16'hfafa;
#10;
address_ina = 210;
address_inb = 211;
data_ina = 16'h23c;
data_inb = 16'h314;
#10;
address_ina = 212;
address_inb = 213;
data_ina = 16'hfb28;
data_inb = 16'hfc8e;
#10;
address_ina = 214;
address_inb = 215;
data_ina = 16'he;
data_inb = 16'h4cf;
#10;
address_ina = 216;
address_inb = 217;
data_ina = 16'h27b;
data_inb = 16'hff6d;
#10;
address_ina = 218;
address_inb = 219;
data_ina = 16'hfa33;
data_inb = 16'hfebe;
#10;
address_ina = 220;
address_inb = 221;
data_ina = 16'h147;
data_inb = 16'h64a;
#10;
address_ina = 222;
address_inb = 223;
data_ina = 16'h348;
data_inb = 16'h3e2;
#10;
address_ina = 224;
address_inb = 225;
data_ina = 16'he7;
data_inb = 16'hfb54;
#10;
address_ina = 226;
address_inb = 227;
data_ina = 16'h649;
data_inb = 16'h57f;
#10;
address_ina = 228;
address_inb = 229;
data_ina = 16'hfa6e;
data_inb = 16'h209;
#10;
address_ina = 230;
address_inb = 231;
data_ina = 16'h587;
data_inb = 16'h214;
#10;
address_ina = 232;
address_inb = 233;
data_ina = 16'hfe71;
data_inb = 16'hfdfc;
#10;
address_ina = 234;
address_inb = 235;
data_ina = 16'hfb24;
data_inb = 16'hfd7b;
#10;
address_ina = 236;
address_inb = 237;
data_ina = 16'hfdb0;
data_inb = 16'hfe22;
#10;
address_ina = 238;
address_inb = 239;
data_ina = 16'h3c9;
data_inb = 16'hfcd9;
#10;
address_ina = 240;
address_inb = 241;
data_ina = 16'h3d9;
data_inb = 16'h11e;
#10;
address_ina = 242;
address_inb = 243;
data_ina = 16'h440;
data_inb = 16'hfac7;
#10;
address_ina = 244;
address_inb = 245;
data_ina = 16'h66d;
data_inb = 16'hfad0;
#10;
address_ina = 246;
address_inb = 247;
data_ina = 16'hfd31;
data_inb = 16'h371;
#10;
address_ina = 248;
address_inb = 249;
data_ina = 16'hfa51;
data_inb = 16'h382;
#10;
address_ina = 250;
address_inb = 251;
data_ina = 16'h67d;
data_inb = 16'hfc17;
#10;
address_ina = 252;
address_inb = 253;
data_ina = 16'h4f7;
data_inb = 16'hfb;
#10;
address_ina = 254;
address_inb = 255;
data_ina = 16'h4e2;
data_inb = 16'h659;
#10;
        wait(init_done);
        #30
        we = 0;
        // Start processing
         
		  #38000

        start = 0;



//        wait (wr_req);
//		  wait (!wr_req);
//		   rd_req = 1;
		  wait(done);
		  #20000
rd_req = 1;
        #70 
		  start = 1;
		 #80 
wait(rd_empty)
rd_req = 0;

$display("Finished the NTT test Number %d",test_num);
////Begin test number #84//////////////
rst = 1;

//#1000
start = 1;
mode = 1; //NTT 0 // INTT 1

// Reset for a few clock cycles

#1000

rst = 0;
test_num = test_num + 1;
#1000
we = 1;
address_ina = 0;
address_inb = 1;
data_ina = 16'hf9e7;
data_inb = 16'h3a3;
#10;
address_ina = 2;
address_inb = 3;
data_ina = 16'hfab1;
data_inb = 16'h372;
#10;
address_ina = 4;
address_inb = 5;
data_ina = 16'hfa0f;
data_inb = 16'hfd51;
#10;
address_ina = 6;
address_inb = 7;
data_ina = 16'h2d6;
data_inb = 16'hf986;
#10;
address_ina = 8;
address_inb = 9;
data_ina = 16'hfadb;
data_inb = 16'h63d;
#10;
address_ina = 10;
address_inb = 11;
data_ina = 16'hff3a;
data_inb = 16'hfc91;
#10;
address_ina = 12;
address_inb = 13;
data_ina = 16'h1a4;
data_inb = 16'hfca8;
#10;
address_ina = 14;
address_inb = 15;
data_ina = 16'hfb30;
data_inb = 16'hfc1c;
#10;
address_ina = 16;
address_inb = 17;
data_ina = 16'hfd51;
data_inb = 16'hfae2;
#10;
address_ina = 18;
address_inb = 19;
data_ina = 16'hff47;
data_inb = 16'h2db;
#10;
address_ina = 20;
address_inb = 21;
data_ina = 16'h85;
data_inb = 16'hfa02;
#10;
address_ina = 22;
address_inb = 23;
data_ina = 16'h135;
data_inb = 16'hfb3f;
#10;
address_ina = 24;
address_inb = 25;
data_ina = 16'h366;
data_inb = 16'hfcb7;
#10;
address_ina = 26;
address_inb = 27;
data_ina = 16'hfdd6;
data_inb = 16'hfe60;
#10;
address_ina = 28;
address_inb = 29;
data_ina = 16'hfda9;
data_inb = 16'hff51;
#10;
address_ina = 30;
address_inb = 31;
data_ina = 16'hfd02;
data_inb = 16'hfbfe;
#10;
address_ina = 32;
address_inb = 33;
data_ina = 16'hfa09;
data_inb = 16'h5b7;
#10;
address_ina = 34;
address_inb = 35;
data_ina = 16'hfcfb;
data_inb = 16'h619;
#10;
address_ina = 36;
address_inb = 37;
data_ina = 16'h549;
data_inb = 16'h1a9;
#10;
address_ina = 38;
address_inb = 39;
data_ina = 16'h651;
data_inb = 16'h249;
#10;
address_ina = 40;
address_inb = 41;
data_ina = 16'hfb21;
data_inb = 16'h2d1;
#10;
address_ina = 42;
address_inb = 43;
data_ina = 16'hfe81;
data_inb = 16'hfcce;
#10;
address_ina = 44;
address_inb = 45;
data_ina = 16'hfbe6;
data_inb = 16'hf9ff;
#10;
address_ina = 46;
address_inb = 47;
data_ina = 16'h372;
data_inb = 16'h1d2;
#10;
address_ina = 48;
address_inb = 49;
data_ina = 16'hc2;
data_inb = 16'hfb30;
#10;
address_ina = 50;
address_inb = 51;
data_ina = 16'hfe3a;
data_inb = 16'h3e6;
#10;
address_ina = 52;
address_inb = 53;
data_ina = 16'h3f;
data_inb = 16'hf9b7;
#10;
address_ina = 54;
address_inb = 55;
data_ina = 16'hfd63;
data_inb = 16'h550;
#10;
address_ina = 56;
address_inb = 57;
data_ina = 16'hfe4f;
data_inb = 16'h1c1;
#10;
address_ina = 58;
address_inb = 59;
data_ina = 16'hff9c;
data_inb = 16'hfe14;
#10;
address_ina = 60;
address_inb = 61;
data_ina = 16'h87;
data_inb = 16'h15b;
#10;
address_ina = 62;
address_inb = 63;
data_ina = 16'hfab2;
data_inb = 16'had;
#10;
address_ina = 64;
address_inb = 65;
data_ina = 16'hfc49;
data_inb = 16'h3c;
#10;
address_ina = 66;
address_inb = 67;
data_ina = 16'hf9d4;
data_inb = 16'h55f;
#10;
address_ina = 68;
address_inb = 69;
data_ina = 16'hfe9f;
data_inb = 16'hff86;
#10;
address_ina = 70;
address_inb = 71;
data_ina = 16'hfb50;
data_inb = 16'h55f;
#10;
address_ina = 72;
address_inb = 73;
data_ina = 16'hfe18;
data_inb = 16'h1e7;
#10;
address_ina = 74;
address_inb = 75;
data_ina = 16'hfaa7;
data_inb = 16'hfcff;
#10;
address_ina = 76;
address_inb = 77;
data_ina = 16'h3f4;
data_inb = 16'h350;
#10;
address_ina = 78;
address_inb = 79;
data_ina = 16'hfbab;
data_inb = 16'hfa77;
#10;
address_ina = 80;
address_inb = 81;
data_ina = 16'h528;
data_inb = 16'h47f;
#10;
address_ina = 82;
address_inb = 83;
data_ina = 16'h429;
data_inb = 16'hfb61;
#10;
address_ina = 84;
address_inb = 85;
data_ina = 16'hfab6;
data_inb = 16'ha5;
#10;
address_ina = 86;
address_inb = 87;
data_ina = 16'h4ca;
data_inb = 16'hfdc1;
#10;
address_ina = 88;
address_inb = 89;
data_ina = 16'h54a;
data_inb = 16'h4ba;
#10;
address_ina = 90;
address_inb = 91;
data_ina = 16'hfb9e;
data_inb = 16'hfce4;
#10;
address_ina = 92;
address_inb = 93;
data_ina = 16'hff9e;
data_inb = 16'hfc5a;
#10;
address_ina = 94;
address_inb = 95;
data_ina = 16'hfd2a;
data_inb = 16'hfc89;
#10;
address_ina = 96;
address_inb = 97;
data_ina = 16'h57d;
data_inb = 16'hfd1b;
#10;
address_ina = 98;
address_inb = 99;
data_ina = 16'hffb7;
data_inb = 16'h630;
#10;
address_ina = 100;
address_inb = 101;
data_ina = 16'hfe50;
data_inb = 16'h93;
#10;
address_ina = 102;
address_inb = 103;
data_ina = 16'h413;
data_inb = 16'h66c;
#10;
address_ina = 104;
address_inb = 105;
data_ina = 16'hfd68;
data_inb = 16'h16c;
#10;
address_ina = 106;
address_inb = 107;
data_ina = 16'hfe65;
data_inb = 16'h56a;
#10;
address_ina = 108;
address_inb = 109;
data_ina = 16'h2cb;
data_inb = 16'h5f1;
#10;
address_ina = 110;
address_inb = 111;
data_ina = 16'hfd60;
data_inb = 16'h45b;
#10;
address_ina = 112;
address_inb = 113;
data_ina = 16'h660;
data_inb = 16'h51d;
#10;
address_ina = 114;
address_inb = 115;
data_ina = 16'h30b;
data_inb = 16'h211;
#10;
address_ina = 116;
address_inb = 117;
data_ina = 16'hf9d0;
data_inb = 16'h245;
#10;
address_ina = 118;
address_inb = 119;
data_ina = 16'hfc11;
data_inb = 16'h3c9;
#10;
address_ina = 120;
address_inb = 121;
data_ina = 16'hfd88;
data_inb = 16'hfe3d;
#10;
address_ina = 122;
address_inb = 123;
data_ina = 16'h2f9;
data_inb = 16'hfb13;
#10;
address_ina = 124;
address_inb = 125;
data_ina = 16'hfef5;
data_inb = 16'hfc4f;
#10;
address_ina = 126;
address_inb = 127;
data_ina = 16'hffbc;
data_inb = 16'hfb46;
#10;
address_ina = 128;
address_inb = 129;
data_ina = 16'h50f;
data_inb = 16'hde;
#10;
address_ina = 130;
address_inb = 131;
data_ina = 16'hfecc;
data_inb = 16'hfcba;
#10;
address_ina = 132;
address_inb = 133;
data_ina = 16'h41a;
data_inb = 16'hfc3d;
#10;
address_ina = 134;
address_inb = 135;
data_ina = 16'h672;
data_inb = 16'h25e;
#10;
address_ina = 136;
address_inb = 137;
data_ina = 16'h440;
data_inb = 16'h1f9;
#10;
address_ina = 138;
address_inb = 139;
data_ina = 16'h246;
data_inb = 16'h105;
#10;
address_ina = 140;
address_inb = 141;
data_ina = 16'hfb38;
data_inb = 16'h23d;
#10;
address_ina = 142;
address_inb = 143;
data_ina = 16'h174;
data_inb = 16'hfb39;
#10;
address_ina = 144;
address_inb = 145;
data_ina = 16'h615;
data_inb = 16'hfbc1;
#10;
address_ina = 146;
address_inb = 147;
data_ina = 16'h4c2;
data_inb = 16'hfe17;
#10;
address_ina = 148;
address_inb = 149;
data_ina = 16'hfcf6;
data_inb = 16'hfa85;
#10;
address_ina = 150;
address_inb = 151;
data_ina = 16'h352;
data_inb = 16'hfb72;
#10;
address_ina = 152;
address_inb = 153;
data_ina = 16'h677;
data_inb = 16'hca;
#10;
address_ina = 154;
address_inb = 155;
data_ina = 16'h58e;
data_inb = 16'h31d;
#10;
address_ina = 156;
address_inb = 157;
data_ina = 16'h35f;
data_inb = 16'hff1f;
#10;
address_ina = 158;
address_inb = 159;
data_ina = 16'hfd82;
data_inb = 16'hfb27;
#10;
address_ina = 160;
address_inb = 161;
data_ina = 16'hff87;
data_inb = 16'h586;
#10;
address_ina = 162;
address_inb = 163;
data_ina = 16'hfa57;
data_inb = 16'h2cf;
#10;
address_ina = 164;
address_inb = 165;
data_ina = 16'hffc6;
data_inb = 16'hff74;
#10;
address_ina = 166;
address_inb = 167;
data_ina = 16'hfe59;
data_inb = 16'hfb58;
#10;
address_ina = 168;
address_inb = 169;
data_ina = 16'hfc7d;
data_inb = 16'h119;
#10;
address_ina = 170;
address_inb = 171;
data_ina = 16'hfc3d;
data_inb = 16'h1a;
#10;
address_ina = 172;
address_inb = 173;
data_ina = 16'h232;
data_inb = 16'hc8;
#10;
address_ina = 174;
address_inb = 175;
data_ina = 16'hf99a;
data_inb = 16'hf983;
#10;
address_ina = 176;
address_inb = 177;
data_ina = 16'hfcbd;
data_inb = 16'h4d6;
#10;
address_ina = 178;
address_inb = 179;
data_ina = 16'hfe3d;
data_inb = 16'h1e;
#10;
address_ina = 180;
address_inb = 181;
data_ina = 16'h3f8;
data_inb = 16'hfe35;
#10;
address_ina = 182;
address_inb = 183;
data_ina = 16'h75;
data_inb = 16'hfba6;
#10;
address_ina = 184;
address_inb = 185;
data_ina = 16'hfff5;
data_inb = 16'hfdb3;
#10;
address_ina = 186;
address_inb = 187;
data_ina = 16'h1fc;
data_inb = 16'h43a;
#10;
address_ina = 188;
address_inb = 189;
data_ina = 16'hfced;
data_inb = 16'h28e;
#10;
address_ina = 190;
address_inb = 191;
data_ina = 16'h50a;
data_inb = 16'hf9;
#10;
address_ina = 192;
address_inb = 193;
data_ina = 16'hfc28;
data_inb = 16'hfe5d;
#10;
address_ina = 194;
address_inb = 195;
data_ina = 16'h40c;
data_inb = 16'h62d;
#10;
address_ina = 196;
address_inb = 197;
data_ina = 16'h128;
data_inb = 16'hfd25;
#10;
address_ina = 198;
address_inb = 199;
data_ina = 16'h29b;
data_inb = 16'h88;
#10;
address_ina = 200;
address_inb = 201;
data_ina = 16'h35d;
data_inb = 16'h660;
#10;
address_ina = 202;
address_inb = 203;
data_ina = 16'hf9d3;
data_inb = 16'h409;
#10;
address_ina = 204;
address_inb = 205;
data_ina = 16'hfb3a;
data_inb = 16'h160;
#10;
address_ina = 206;
address_inb = 207;
data_ina = 16'h21b;
data_inb = 16'h112;
#10;
address_ina = 208;
address_inb = 209;
data_ina = 16'hfede;
data_inb = 16'he6;
#10;
address_ina = 210;
address_inb = 211;
data_ina = 16'hfda2;
data_inb = 16'hff3b;
#10;
address_ina = 212;
address_inb = 213;
data_ina = 16'hfd67;
data_inb = 16'h3c1;
#10;
address_ina = 214;
address_inb = 215;
data_ina = 16'hfe34;
data_inb = 16'hfa8c;
#10;
address_ina = 216;
address_inb = 217;
data_ina = 16'hfbd9;
data_inb = 16'hfa0c;
#10;
address_ina = 218;
address_inb = 219;
data_ina = 16'hfe0c;
data_inb = 16'hff1f;
#10;
address_ina = 220;
address_inb = 221;
data_ina = 16'hffed;
data_inb = 16'h225;
#10;
address_ina = 222;
address_inb = 223;
data_ina = 16'h483;
data_inb = 16'h320;
#10;
address_ina = 224;
address_inb = 225;
data_ina = 16'hfd55;
data_inb = 16'hfc9c;
#10;
address_ina = 226;
address_inb = 227;
data_ina = 16'h43e;
data_inb = 16'h243;
#10;
address_ina = 228;
address_inb = 229;
data_ina = 16'hfc68;
data_inb = 16'h618;
#10;
address_ina = 230;
address_inb = 231;
data_ina = 16'hfa3e;
data_inb = 16'h5a9;
#10;
address_ina = 232;
address_inb = 233;
data_ina = 16'h360;
data_inb = 16'hfa6d;
#10;
address_ina = 234;
address_inb = 235;
data_ina = 16'h3fa;
data_inb = 16'h166;
#10;
address_ina = 236;
address_inb = 237;
data_ina = 16'h652;
data_inb = 16'hfc59;
#10;
address_ina = 238;
address_inb = 239;
data_ina = 16'hff08;
data_inb = 16'hf99f;
#10;
address_ina = 240;
address_inb = 241;
data_ina = 16'hfe18;
data_inb = 16'h1bf;
#10;
address_ina = 242;
address_inb = 243;
data_ina = 16'h3d7;
data_inb = 16'hfb38;
#10;
address_ina = 244;
address_inb = 245;
data_ina = 16'hfe29;
data_inb = 16'hff0f;
#10;
address_ina = 246;
address_inb = 247;
data_ina = 16'hfccc;
data_inb = 16'hfd0e;
#10;
address_ina = 248;
address_inb = 249;
data_ina = 16'hdf;
data_inb = 16'hb4;
#10;
address_ina = 250;
address_inb = 251;
data_ina = 16'hfc6f;
data_inb = 16'h60b;
#10;
address_ina = 252;
address_inb = 253;
data_ina = 16'h25e;
data_inb = 16'hfbc6;
#10;
address_ina = 254;
address_inb = 255;
data_ina = 16'hd3;
data_inb = 16'hfff5;
#10;
        wait(init_done);
        #30
        we = 0;
        // Start processing
         
		  #38000

        start = 0;



//        wait (wr_req);
//		  wait (!wr_req);
//		   rd_req = 1;
		  wait(done);
		  #20000
rd_req = 1;
        #70 
		  start = 1;
		 #80 
wait(rd_empty)
rd_req = 0;

$display("Finished the NTT test Number %d",test_num);
////Begin test number #85//////////////
rst = 1;

//#1000
start = 1;
mode = 0; //NTT 0 // INTT 1

// Reset for a few clock cycles

#1000

rst = 0;
test_num = test_num + 1;
#1000
we = 1;
address_ina = 0;
address_inb = 1;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 2;
address_inb = 3;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 4;
address_inb = 5;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 6;
address_inb = 7;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 8;
address_inb = 9;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 10;
address_inb = 11;
data_ina = 16'h2;
data_inb = 16'h2;
#10;
address_ina = 12;
address_inb = 13;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 14;
address_inb = 15;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 16;
address_inb = 17;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 18;
address_inb = 19;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 20;
address_inb = 21;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 22;
address_inb = 23;
data_ina = 16'hfffe;
data_inb = 16'hffff;
#10;
address_ina = 24;
address_inb = 25;
data_ina = 16'h3;
data_inb = 16'h0;
#10;
address_ina = 26;
address_inb = 27;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 28;
address_inb = 29;
data_ina = 16'h0;
data_inb = 16'h2;
#10;
address_ina = 30;
address_inb = 31;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 32;
address_inb = 33;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 34;
address_inb = 35;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 36;
address_inb = 37;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 38;
address_inb = 39;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 40;
address_inb = 41;
data_ina = 16'h3;
data_inb = 16'h0;
#10;
address_ina = 42;
address_inb = 43;
data_ina = 16'h1;
data_inb = 16'hfffe;
#10;
address_ina = 44;
address_inb = 45;
data_ina = 16'h0;
data_inb = 16'h2;
#10;
address_ina = 46;
address_inb = 47;
data_ina = 16'h2;
data_inb = 16'hffff;
#10;
address_ina = 48;
address_inb = 49;
data_ina = 16'hfffe;
data_inb = 16'h1;
#10;
address_ina = 50;
address_inb = 51;
data_ina = 16'h0;
data_inb = 16'h2;
#10;
address_ina = 52;
address_inb = 53;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 54;
address_inb = 55;
data_ina = 16'hfffe;
data_inb = 16'h2;
#10;
address_ina = 56;
address_inb = 57;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 58;
address_inb = 59;
data_ina = 16'h2;
data_inb = 16'h3;
#10;
address_ina = 60;
address_inb = 61;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 62;
address_inb = 63;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 64;
address_inb = 65;
data_ina = 16'h1;
data_inb = 16'h2;
#10;
address_ina = 66;
address_inb = 67;
data_ina = 16'h2;
data_inb = 16'h0;
#10;
address_ina = 68;
address_inb = 69;
data_ina = 16'hfffd;
data_inb = 16'h1;
#10;
address_ina = 70;
address_inb = 71;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 72;
address_inb = 73;
data_ina = 16'hfffe;
data_inb = 16'h1;
#10;
address_ina = 74;
address_inb = 75;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 76;
address_inb = 77;
data_ina = 16'hfffe;
data_inb = 16'hffff;
#10;
address_ina = 78;
address_inb = 79;
data_ina = 16'hffff;
data_inb = 16'h2;
#10;
address_ina = 80;
address_inb = 81;
data_ina = 16'h1;
data_inb = 16'h2;
#10;
address_ina = 82;
address_inb = 83;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 84;
address_inb = 85;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 86;
address_inb = 87;
data_ina = 16'hfffe;
data_inb = 16'h0;
#10;
address_ina = 88;
address_inb = 89;
data_ina = 16'h2;
data_inb = 16'h1;
#10;
address_ina = 90;
address_inb = 91;
data_ina = 16'hfffe;
data_inb = 16'hffff;
#10;
address_ina = 92;
address_inb = 93;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 94;
address_inb = 95;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 96;
address_inb = 97;
data_ina = 16'hfffd;
data_inb = 16'hfffe;
#10;
address_ina = 98;
address_inb = 99;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 100;
address_inb = 101;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 102;
address_inb = 103;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 104;
address_inb = 105;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 106;
address_inb = 107;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 108;
address_inb = 109;
data_ina = 16'h1;
data_inb = 16'hfffd;
#10;
address_ina = 110;
address_inb = 111;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 112;
address_inb = 113;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 114;
address_inb = 115;
data_ina = 16'h1;
data_inb = 16'h2;
#10;
address_ina = 116;
address_inb = 117;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 118;
address_inb = 119;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 120;
address_inb = 121;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 122;
address_inb = 123;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 124;
address_inb = 125;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 126;
address_inb = 127;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 128;
address_inb = 129;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 130;
address_inb = 131;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 132;
address_inb = 133;
data_ina = 16'h1;
data_inb = 16'h2;
#10;
address_ina = 134;
address_inb = 135;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 136;
address_inb = 137;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 138;
address_inb = 139;
data_ina = 16'h0;
data_inb = 16'hfffe;
#10;
address_ina = 140;
address_inb = 141;
data_ina = 16'hfffe;
data_inb = 16'hffff;
#10;
address_ina = 142;
address_inb = 143;
data_ina = 16'h0;
data_inb = 16'h2;
#10;
address_ina = 144;
address_inb = 145;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 146;
address_inb = 147;
data_ina = 16'h2;
data_inb = 16'h1;
#10;
address_ina = 148;
address_inb = 149;
data_ina = 16'hfffe;
data_inb = 16'hffff;
#10;
address_ina = 150;
address_inb = 151;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 152;
address_inb = 153;
data_ina = 16'hffff;
data_inb = 16'hfffe;
#10;
address_ina = 154;
address_inb = 155;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 156;
address_inb = 157;
data_ina = 16'hfffe;
data_inb = 16'h1;
#10;
address_ina = 158;
address_inb = 159;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 160;
address_inb = 161;
data_ina = 16'h2;
data_inb = 16'hffff;
#10;
address_ina = 162;
address_inb = 163;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 164;
address_inb = 165;
data_ina = 16'h2;
data_inb = 16'h0;
#10;
address_ina = 166;
address_inb = 167;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 168;
address_inb = 169;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 170;
address_inb = 171;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 172;
address_inb = 173;
data_ina = 16'h2;
data_inb = 16'h1;
#10;
address_ina = 174;
address_inb = 175;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 176;
address_inb = 177;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 178;
address_inb = 179;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 180;
address_inb = 181;
data_ina = 16'hffff;
data_inb = 16'hfffd;
#10;
address_ina = 182;
address_inb = 183;
data_ina = 16'h1;
data_inb = 16'hfffe;
#10;
address_ina = 184;
address_inb = 185;
data_ina = 16'h0;
data_inb = 16'h2;
#10;
address_ina = 186;
address_inb = 187;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 188;
address_inb = 189;
data_ina = 16'hfffe;
data_inb = 16'hffff;
#10;
address_ina = 190;
address_inb = 191;
data_ina = 16'h1;
data_inb = 16'h2;
#10;
address_ina = 192;
address_inb = 193;
data_ina = 16'hffff;
data_inb = 16'h2;
#10;
address_ina = 194;
address_inb = 195;
data_ina = 16'h2;
data_inb = 16'h0;
#10;
address_ina = 196;
address_inb = 197;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 198;
address_inb = 199;
data_ina = 16'hffff;
data_inb = 16'hfffe;
#10;
address_ina = 200;
address_inb = 201;
data_ina = 16'h1;
data_inb = 16'h2;
#10;
address_ina = 202;
address_inb = 203;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 204;
address_inb = 205;
data_ina = 16'h2;
data_inb = 16'h1;
#10;
address_ina = 206;
address_inb = 207;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 208;
address_inb = 209;
data_ina = 16'h2;
data_inb = 16'hffff;
#10;
address_ina = 210;
address_inb = 211;
data_ina = 16'hffff;
data_inb = 16'hfffe;
#10;
address_ina = 212;
address_inb = 213;
data_ina = 16'h2;
data_inb = 16'h0;
#10;
address_ina = 214;
address_inb = 215;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 216;
address_inb = 217;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 218;
address_inb = 219;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 220;
address_inb = 221;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 222;
address_inb = 223;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 224;
address_inb = 225;
data_ina = 16'h2;
data_inb = 16'h1;
#10;
address_ina = 226;
address_inb = 227;
data_ina = 16'h1;
data_inb = 16'h2;
#10;
address_ina = 228;
address_inb = 229;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 230;
address_inb = 231;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 232;
address_inb = 233;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 234;
address_inb = 235;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 236;
address_inb = 237;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 238;
address_inb = 239;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 240;
address_inb = 241;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 242;
address_inb = 243;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 244;
address_inb = 245;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 246;
address_inb = 247;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 248;
address_inb = 249;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 250;
address_inb = 251;
data_ina = 16'hfffd;
data_inb = 16'h0;
#10;
address_ina = 252;
address_inb = 253;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 254;
address_inb = 255;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
        wait(init_done);
        #30
        we = 0;
        // Start processing
         
		  #38000

        start = 0;



//        wait (wr_req);
//		  wait (!wr_req);
//		   rd_req = 1;
		  wait(done);
		  #20000
rd_req = 1;
        #70 
		  start = 1;
		 #80 
wait(rd_empty)
rd_req = 0;

$display("Finished the NTT test Number %d",test_num);
////Begin test number #86//////////////
rst = 1;

//#1000
start = 1;
mode = 0; //NTT 0 // INTT 1

// Reset for a few clock cycles

#1000

rst = 0;
test_num = test_num + 1;
#1000
we = 1;
address_ina = 0;
address_inb = 1;
data_ina = 16'h1;
data_inb = 16'h2;
#10;
address_ina = 2;
address_inb = 3;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 4;
address_inb = 5;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 6;
address_inb = 7;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 8;
address_inb = 9;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 10;
address_inb = 11;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 12;
address_inb = 13;
data_ina = 16'hfffe;
data_inb = 16'h1;
#10;
address_ina = 14;
address_inb = 15;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 16;
address_inb = 17;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 18;
address_inb = 19;
data_ina = 16'h0;
data_inb = 16'hfffe;
#10;
address_ina = 20;
address_inb = 21;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 22;
address_inb = 23;
data_ina = 16'h0;
data_inb = 16'hfffe;
#10;
address_ina = 24;
address_inb = 25;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 26;
address_inb = 27;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 28;
address_inb = 29;
data_ina = 16'h1;
data_inb = 16'h2;
#10;
address_ina = 30;
address_inb = 31;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 32;
address_inb = 33;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 34;
address_inb = 35;
data_ina = 16'hfffe;
data_inb = 16'h0;
#10;
address_ina = 36;
address_inb = 37;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 38;
address_inb = 39;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 40;
address_inb = 41;
data_ina = 16'hffff;
data_inb = 16'h2;
#10;
address_ina = 42;
address_inb = 43;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 44;
address_inb = 45;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 46;
address_inb = 47;
data_ina = 16'h0;
data_inb = 16'hfffe;
#10;
address_ina = 48;
address_inb = 49;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 50;
address_inb = 51;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 52;
address_inb = 53;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 54;
address_inb = 55;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 56;
address_inb = 57;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 58;
address_inb = 59;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 60;
address_inb = 61;
data_ina = 16'h0;
data_inb = 16'hfffe;
#10;
address_ina = 62;
address_inb = 63;
data_ina = 16'h0;
data_inb = 16'h3;
#10;
address_ina = 64;
address_inb = 65;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 66;
address_inb = 67;
data_ina = 16'hffff;
data_inb = 16'hfffe;
#10;
address_ina = 68;
address_inb = 69;
data_ina = 16'hffff;
data_inb = 16'h2;
#10;
address_ina = 70;
address_inb = 71;
data_ina = 16'h2;
data_inb = 16'hffff;
#10;
address_ina = 72;
address_inb = 73;
data_ina = 16'h2;
data_inb = 16'h1;
#10;
address_ina = 74;
address_inb = 75;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 76;
address_inb = 77;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 78;
address_inb = 79;
data_ina = 16'hffff;
data_inb = 16'hfffd;
#10;
address_ina = 80;
address_inb = 81;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 82;
address_inb = 83;
data_ina = 16'h2;
data_inb = 16'h0;
#10;
address_ina = 84;
address_inb = 85;
data_ina = 16'h0;
data_inb = 16'hfffe;
#10;
address_ina = 86;
address_inb = 87;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 88;
address_inb = 89;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 90;
address_inb = 91;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 92;
address_inb = 93;
data_ina = 16'h2;
data_inb = 16'h1;
#10;
address_ina = 94;
address_inb = 95;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 96;
address_inb = 97;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 98;
address_inb = 99;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 100;
address_inb = 101;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 102;
address_inb = 103;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 104;
address_inb = 105;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 106;
address_inb = 107;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 108;
address_inb = 109;
data_ina = 16'hffff;
data_inb = 16'hfffd;
#10;
address_ina = 110;
address_inb = 111;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 112;
address_inb = 113;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 114;
address_inb = 115;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 116;
address_inb = 117;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 118;
address_inb = 119;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 120;
address_inb = 121;
data_ina = 16'h1;
data_inb = 16'h2;
#10;
address_ina = 122;
address_inb = 123;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 124;
address_inb = 125;
data_ina = 16'h0;
data_inb = 16'h2;
#10;
address_ina = 126;
address_inb = 127;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 128;
address_inb = 129;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 130;
address_inb = 131;
data_ina = 16'h2;
data_inb = 16'hfffd;
#10;
address_ina = 132;
address_inb = 133;
data_ina = 16'h3;
data_inb = 16'hffff;
#10;
address_ina = 134;
address_inb = 135;
data_ina = 16'hffff;
data_inb = 16'hfffd;
#10;
address_ina = 136;
address_inb = 137;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 138;
address_inb = 139;
data_ina = 16'h2;
data_inb = 16'hffff;
#10;
address_ina = 140;
address_inb = 141;
data_ina = 16'h1;
data_inb = 16'h2;
#10;
address_ina = 142;
address_inb = 143;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 144;
address_inb = 145;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 146;
address_inb = 147;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 148;
address_inb = 149;
data_ina = 16'h0;
data_inb = 16'hfffd;
#10;
address_ina = 150;
address_inb = 151;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 152;
address_inb = 153;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 154;
address_inb = 155;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 156;
address_inb = 157;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 158;
address_inb = 159;
data_ina = 16'hfffd;
data_inb = 16'h1;
#10;
address_ina = 160;
address_inb = 161;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 162;
address_inb = 163;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 164;
address_inb = 165;
data_ina = 16'h0;
data_inb = 16'h2;
#10;
address_ina = 166;
address_inb = 167;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 168;
address_inb = 169;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 170;
address_inb = 171;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 172;
address_inb = 173;
data_ina = 16'hfffe;
data_inb = 16'hffff;
#10;
address_ina = 174;
address_inb = 175;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 176;
address_inb = 177;
data_ina = 16'h1;
data_inb = 16'h2;
#10;
address_ina = 178;
address_inb = 179;
data_ina = 16'h2;
data_inb = 16'h3;
#10;
address_ina = 180;
address_inb = 181;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 182;
address_inb = 183;
data_ina = 16'hfffe;
data_inb = 16'h0;
#10;
address_ina = 184;
address_inb = 185;
data_ina = 16'h2;
data_inb = 16'hffff;
#10;
address_ina = 186;
address_inb = 187;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 188;
address_inb = 189;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 190;
address_inb = 191;
data_ina = 16'hfffe;
data_inb = 16'h1;
#10;
address_ina = 192;
address_inb = 193;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 194;
address_inb = 195;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 196;
address_inb = 197;
data_ina = 16'hfffd;
data_inb = 16'h1;
#10;
address_ina = 198;
address_inb = 199;
data_ina = 16'h1;
data_inb = 16'hfffe;
#10;
address_ina = 200;
address_inb = 201;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 202;
address_inb = 203;
data_ina = 16'hfffe;
data_inb = 16'hffff;
#10;
address_ina = 204;
address_inb = 205;
data_ina = 16'h0;
data_inb = 16'h2;
#10;
address_ina = 206;
address_inb = 207;
data_ina = 16'h2;
data_inb = 16'h1;
#10;
address_ina = 208;
address_inb = 209;
data_ina = 16'h1;
data_inb = 16'hfffe;
#10;
address_ina = 210;
address_inb = 211;
data_ina = 16'hffff;
data_inb = 16'hfffd;
#10;
address_ina = 212;
address_inb = 213;
data_ina = 16'hfffe;
data_inb = 16'h1;
#10;
address_ina = 214;
address_inb = 215;
data_ina = 16'hfffe;
data_inb = 16'h2;
#10;
address_ina = 216;
address_inb = 217;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 218;
address_inb = 219;
data_ina = 16'hfffe;
data_inb = 16'hffff;
#10;
address_ina = 220;
address_inb = 221;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 222;
address_inb = 223;
data_ina = 16'h2;
data_inb = 16'h2;
#10;
address_ina = 224;
address_inb = 225;
data_ina = 16'hfffe;
data_inb = 16'hffff;
#10;
address_ina = 226;
address_inb = 227;
data_ina = 16'hfffe;
data_inb = 16'h1;
#10;
address_ina = 228;
address_inb = 229;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 230;
address_inb = 231;
data_ina = 16'h2;
data_inb = 16'h0;
#10;
address_ina = 232;
address_inb = 233;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 234;
address_inb = 235;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 236;
address_inb = 237;
data_ina = 16'h0;
data_inb = 16'h2;
#10;
address_ina = 238;
address_inb = 239;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 240;
address_inb = 241;
data_ina = 16'h2;
data_inb = 16'hfffe;
#10;
address_ina = 242;
address_inb = 243;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 244;
address_inb = 245;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 246;
address_inb = 247;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 248;
address_inb = 249;
data_ina = 16'h0;
data_inb = 16'h2;
#10;
address_ina = 250;
address_inb = 251;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 252;
address_inb = 253;
data_ina = 16'h2;
data_inb = 16'hffff;
#10;
address_ina = 254;
address_inb = 255;
data_ina = 16'hffff;
data_inb = 16'hfffe;
#10;
        wait(init_done);
        #30
        we = 0;
        // Start processing
         
		  #38000

        start = 0;



//        wait (wr_req);
//		  wait (!wr_req);
//		   rd_req = 1;
		  wait(done);
		  #20000
rd_req = 1;
        #70 
		  start = 1;
		 #80 
wait(rd_empty)
rd_req = 0;

$display("Finished the NTT test Number %d",test_num);
////Begin test number #87//////////////
rst = 1;

//#1000
start = 1;
mode = 0; //NTT 0 // INTT 1

// Reset for a few clock cycles

#1000

rst = 0;
test_num = test_num + 1;
#1000
we = 1;
address_ina = 0;
address_inb = 1;
data_ina = 16'h0;
data_inb = 16'h2;
#10;
address_ina = 2;
address_inb = 3;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 4;
address_inb = 5;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 6;
address_inb = 7;
data_ina = 16'h2;
data_inb = 16'h1;
#10;
address_ina = 8;
address_inb = 9;
data_ina = 16'hffff;
data_inb = 16'hfffe;
#10;
address_ina = 10;
address_inb = 11;
data_ina = 16'h1;
data_inb = 16'hfffe;
#10;
address_ina = 12;
address_inb = 13;
data_ina = 16'h2;
data_inb = 16'hffff;
#10;
address_ina = 14;
address_inb = 15;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 16;
address_inb = 17;
data_ina = 16'h2;
data_inb = 16'h1;
#10;
address_ina = 18;
address_inb = 19;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 20;
address_inb = 21;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 22;
address_inb = 23;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 24;
address_inb = 25;
data_ina = 16'h1;
data_inb = 16'hfffe;
#10;
address_ina = 26;
address_inb = 27;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 28;
address_inb = 29;
data_ina = 16'hffff;
data_inb = 16'h2;
#10;
address_ina = 30;
address_inb = 31;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 32;
address_inb = 33;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 34;
address_inb = 35;
data_ina = 16'hffff;
data_inb = 16'hfffe;
#10;
address_ina = 36;
address_inb = 37;
data_ina = 16'h2;
data_inb = 16'hffff;
#10;
address_ina = 38;
address_inb = 39;
data_ina = 16'h2;
data_inb = 16'hfffe;
#10;
address_ina = 40;
address_inb = 41;
data_ina = 16'hffff;
data_inb = 16'hfffe;
#10;
address_ina = 42;
address_inb = 43;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 44;
address_inb = 45;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 46;
address_inb = 47;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 48;
address_inb = 49;
data_ina = 16'h2;
data_inb = 16'hffff;
#10;
address_ina = 50;
address_inb = 51;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 52;
address_inb = 53;
data_ina = 16'hfffe;
data_inb = 16'h0;
#10;
address_ina = 54;
address_inb = 55;
data_ina = 16'h1;
data_inb = 16'h2;
#10;
address_ina = 56;
address_inb = 57;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 58;
address_inb = 59;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 60;
address_inb = 61;
data_ina = 16'hfffe;
data_inb = 16'h0;
#10;
address_ina = 62;
address_inb = 63;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 64;
address_inb = 65;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 66;
address_inb = 67;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 68;
address_inb = 69;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 70;
address_inb = 71;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 72;
address_inb = 73;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 74;
address_inb = 75;
data_ina = 16'hffff;
data_inb = 16'h3;
#10;
address_ina = 76;
address_inb = 77;
data_ina = 16'hffff;
data_inb = 16'hfffe;
#10;
address_ina = 78;
address_inb = 79;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 80;
address_inb = 81;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 82;
address_inb = 83;
data_ina = 16'h2;
data_inb = 16'h0;
#10;
address_ina = 84;
address_inb = 85;
data_ina = 16'hfffe;
data_inb = 16'h1;
#10;
address_ina = 86;
address_inb = 87;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 88;
address_inb = 89;
data_ina = 16'h0;
data_inb = 16'hfffe;
#10;
address_ina = 90;
address_inb = 91;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 92;
address_inb = 93;
data_ina = 16'hffff;
data_inb = 16'h2;
#10;
address_ina = 94;
address_inb = 95;
data_ina = 16'h0;
data_inb = 16'h3;
#10;
address_ina = 96;
address_inb = 97;
data_ina = 16'h0;
data_inb = 16'h2;
#10;
address_ina = 98;
address_inb = 99;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 100;
address_inb = 101;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 102;
address_inb = 103;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 104;
address_inb = 105;
data_ina = 16'h2;
data_inb = 16'hfffe;
#10;
address_ina = 106;
address_inb = 107;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 108;
address_inb = 109;
data_ina = 16'hffff;
data_inb = 16'h2;
#10;
address_ina = 110;
address_inb = 111;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 112;
address_inb = 113;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 114;
address_inb = 115;
data_ina = 16'hfffe;
data_inb = 16'h0;
#10;
address_ina = 116;
address_inb = 117;
data_ina = 16'h1;
data_inb = 16'hfffe;
#10;
address_ina = 118;
address_inb = 119;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 120;
address_inb = 121;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 122;
address_inb = 123;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 124;
address_inb = 125;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 126;
address_inb = 127;
data_ina = 16'h0;
data_inb = 16'h2;
#10;
address_ina = 128;
address_inb = 129;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 130;
address_inb = 131;
data_ina = 16'h2;
data_inb = 16'h2;
#10;
address_ina = 132;
address_inb = 133;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 134;
address_inb = 135;
data_ina = 16'hfffe;
data_inb = 16'h0;
#10;
address_ina = 136;
address_inb = 137;
data_ina = 16'h2;
data_inb = 16'h0;
#10;
address_ina = 138;
address_inb = 139;
data_ina = 16'h2;
data_inb = 16'hfffd;
#10;
address_ina = 140;
address_inb = 141;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 142;
address_inb = 143;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 144;
address_inb = 145;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 146;
address_inb = 147;
data_ina = 16'h2;
data_inb = 16'hffff;
#10;
address_ina = 148;
address_inb = 149;
data_ina = 16'h1;
data_inb = 16'h2;
#10;
address_ina = 150;
address_inb = 151;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 152;
address_inb = 153;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 154;
address_inb = 155;
data_ina = 16'h1;
data_inb = 16'hfffe;
#10;
address_ina = 156;
address_inb = 157;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 158;
address_inb = 159;
data_ina = 16'hfffe;
data_inb = 16'h0;
#10;
address_ina = 160;
address_inb = 161;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 162;
address_inb = 163;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 164;
address_inb = 165;
data_ina = 16'hfffe;
data_inb = 16'h1;
#10;
address_ina = 166;
address_inb = 167;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 168;
address_inb = 169;
data_ina = 16'h2;
data_inb = 16'hffff;
#10;
address_ina = 170;
address_inb = 171;
data_ina = 16'hfffe;
data_inb = 16'hffff;
#10;
address_ina = 172;
address_inb = 173;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 174;
address_inb = 175;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 176;
address_inb = 177;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 178;
address_inb = 179;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 180;
address_inb = 181;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 182;
address_inb = 183;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 184;
address_inb = 185;
data_ina = 16'h0;
data_inb = 16'h2;
#10;
address_ina = 186;
address_inb = 187;
data_ina = 16'h1;
data_inb = 16'h2;
#10;
address_ina = 188;
address_inb = 189;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 190;
address_inb = 191;
data_ina = 16'hffff;
data_inb = 16'hfffd;
#10;
address_ina = 192;
address_inb = 193;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 194;
address_inb = 195;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 196;
address_inb = 197;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 198;
address_inb = 199;
data_ina = 16'h2;
data_inb = 16'hffff;
#10;
address_ina = 200;
address_inb = 201;
data_ina = 16'hfffe;
data_inb = 16'h0;
#10;
address_ina = 202;
address_inb = 203;
data_ina = 16'hfffd;
data_inb = 16'h0;
#10;
address_ina = 204;
address_inb = 205;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 206;
address_inb = 207;
data_ina = 16'hfffe;
data_inb = 16'hffff;
#10;
address_ina = 208;
address_inb = 209;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 210;
address_inb = 211;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 212;
address_inb = 213;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 214;
address_inb = 215;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 216;
address_inb = 217;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 218;
address_inb = 219;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 220;
address_inb = 221;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 222;
address_inb = 223;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 224;
address_inb = 225;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 226;
address_inb = 227;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 228;
address_inb = 229;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 230;
address_inb = 231;
data_ina = 16'hfffe;
data_inb = 16'hffff;
#10;
address_ina = 232;
address_inb = 233;
data_ina = 16'hfffe;
data_inb = 16'h1;
#10;
address_ina = 234;
address_inb = 235;
data_ina = 16'hfffe;
data_inb = 16'h1;
#10;
address_ina = 236;
address_inb = 237;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 238;
address_inb = 239;
data_ina = 16'h0;
data_inb = 16'hfffe;
#10;
address_ina = 240;
address_inb = 241;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 242;
address_inb = 243;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 244;
address_inb = 245;
data_ina = 16'hffff;
data_inb = 16'h3;
#10;
address_ina = 246;
address_inb = 247;
data_ina = 16'h3;
data_inb = 16'hfffe;
#10;
address_ina = 248;
address_inb = 249;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 250;
address_inb = 251;
data_ina = 16'h0;
data_inb = 16'h2;
#10;
address_ina = 252;
address_inb = 253;
data_ina = 16'h2;
data_inb = 16'h1;
#10;
address_ina = 254;
address_inb = 255;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
        wait(init_done);
        #30
        we = 0;
        // Start processing
         
		  #38000

        start = 0;



//        wait (wr_req);
//		  wait (!wr_req);
//		   rd_req = 1;
		  wait(done);
		  #20000
rd_req = 1;
        #70 
		  start = 1;
		 #80 
wait(rd_empty)
rd_req = 0;

$display("Finished the NTT test Number %d",test_num);
////Begin test number #88//////////////
rst = 1;

//#1000
start = 1;
mode = 0; //NTT 0 // INTT 1

// Reset for a few clock cycles

#1000

rst = 0;
test_num = test_num + 1;
#1000
we = 1;
address_ina = 0;
address_inb = 1;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 2;
address_inb = 3;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 4;
address_inb = 5;
data_ina = 16'h1;
data_inb = 16'hfffe;
#10;
address_ina = 6;
address_inb = 7;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 8;
address_inb = 9;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 10;
address_inb = 11;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 12;
address_inb = 13;
data_ina = 16'h2;
data_inb = 16'h1;
#10;
address_ina = 14;
address_inb = 15;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 16;
address_inb = 17;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 18;
address_inb = 19;
data_ina = 16'h3;
data_inb = 16'h0;
#10;
address_ina = 20;
address_inb = 21;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 22;
address_inb = 23;
data_ina = 16'h1;
data_inb = 16'h3;
#10;
address_ina = 24;
address_inb = 25;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 26;
address_inb = 27;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 28;
address_inb = 29;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 30;
address_inb = 31;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 32;
address_inb = 33;
data_ina = 16'hffff;
data_inb = 16'h2;
#10;
address_ina = 34;
address_inb = 35;
data_ina = 16'hffff;
data_inb = 16'h2;
#10;
address_ina = 36;
address_inb = 37;
data_ina = 16'h0;
data_inb = 16'hfffe;
#10;
address_ina = 38;
address_inb = 39;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 40;
address_inb = 41;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 42;
address_inb = 43;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 44;
address_inb = 45;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 46;
address_inb = 47;
data_ina = 16'hffff;
data_inb = 16'h2;
#10;
address_ina = 48;
address_inb = 49;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 50;
address_inb = 51;
data_ina = 16'h1;
data_inb = 16'hfffe;
#10;
address_ina = 52;
address_inb = 53;
data_ina = 16'h1;
data_inb = 16'h2;
#10;
address_ina = 54;
address_inb = 55;
data_ina = 16'h1;
data_inb = 16'h2;
#10;
address_ina = 56;
address_inb = 57;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 58;
address_inb = 59;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 60;
address_inb = 61;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 62;
address_inb = 63;
data_ina = 16'hfffe;
data_inb = 16'hfffd;
#10;
address_ina = 64;
address_inb = 65;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 66;
address_inb = 67;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 68;
address_inb = 69;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 70;
address_inb = 71;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 72;
address_inb = 73;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 74;
address_inb = 75;
data_ina = 16'h2;
data_inb = 16'hffff;
#10;
address_ina = 76;
address_inb = 77;
data_ina = 16'h3;
data_inb = 16'h0;
#10;
address_ina = 78;
address_inb = 79;
data_ina = 16'h2;
data_inb = 16'hffff;
#10;
address_ina = 80;
address_inb = 81;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 82;
address_inb = 83;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 84;
address_inb = 85;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 86;
address_inb = 87;
data_ina = 16'hfffe;
data_inb = 16'h1;
#10;
address_ina = 88;
address_inb = 89;
data_ina = 16'hfffe;
data_inb = 16'h0;
#10;
address_ina = 90;
address_inb = 91;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 92;
address_inb = 93;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 94;
address_inb = 95;
data_ina = 16'h2;
data_inb = 16'h2;
#10;
address_ina = 96;
address_inb = 97;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 98;
address_inb = 99;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 100;
address_inb = 101;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 102;
address_inb = 103;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 104;
address_inb = 105;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 106;
address_inb = 107;
data_ina = 16'hfffd;
data_inb = 16'h1;
#10;
address_ina = 108;
address_inb = 109;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 110;
address_inb = 111;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 112;
address_inb = 113;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 114;
address_inb = 115;
data_ina = 16'h0;
data_inb = 16'hfffe;
#10;
address_ina = 116;
address_inb = 117;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 118;
address_inb = 119;
data_ina = 16'h2;
data_inb = 16'hffff;
#10;
address_ina = 120;
address_inb = 121;
data_ina = 16'hfffe;
data_inb = 16'hffff;
#10;
address_ina = 122;
address_inb = 123;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 124;
address_inb = 125;
data_ina = 16'h2;
data_inb = 16'h1;
#10;
address_ina = 126;
address_inb = 127;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 128;
address_inb = 129;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 130;
address_inb = 131;
data_ina = 16'h1;
data_inb = 16'h3;
#10;
address_ina = 132;
address_inb = 133;
data_ina = 16'h2;
data_inb = 16'h0;
#10;
address_ina = 134;
address_inb = 135;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 136;
address_inb = 137;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 138;
address_inb = 139;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 140;
address_inb = 141;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 142;
address_inb = 143;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 144;
address_inb = 145;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 146;
address_inb = 147;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 148;
address_inb = 149;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 150;
address_inb = 151;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 152;
address_inb = 153;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 154;
address_inb = 155;
data_ina = 16'hfffd;
data_inb = 16'h0;
#10;
address_ina = 156;
address_inb = 157;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 158;
address_inb = 159;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 160;
address_inb = 161;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 162;
address_inb = 163;
data_ina = 16'h0;
data_inb = 16'h2;
#10;
address_ina = 164;
address_inb = 165;
data_ina = 16'h1;
data_inb = 16'hfffe;
#10;
address_ina = 166;
address_inb = 167;
data_ina = 16'h3;
data_inb = 16'h0;
#10;
address_ina = 168;
address_inb = 169;
data_ina = 16'hfffe;
data_inb = 16'hfffe;
#10;
address_ina = 170;
address_inb = 171;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 172;
address_inb = 173;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 174;
address_inb = 175;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 176;
address_inb = 177;
data_ina = 16'hfffe;
data_inb = 16'h0;
#10;
address_ina = 178;
address_inb = 179;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 180;
address_inb = 181;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 182;
address_inb = 183;
data_ina = 16'h1;
data_inb = 16'hfffe;
#10;
address_ina = 184;
address_inb = 185;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 186;
address_inb = 187;
data_ina = 16'hffff;
data_inb = 16'hfffe;
#10;
address_ina = 188;
address_inb = 189;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 190;
address_inb = 191;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 192;
address_inb = 193;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 194;
address_inb = 195;
data_ina = 16'hffff;
data_inb = 16'h2;
#10;
address_ina = 196;
address_inb = 197;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 198;
address_inb = 199;
data_ina = 16'h0;
data_inb = 16'h2;
#10;
address_ina = 200;
address_inb = 201;
data_ina = 16'hffff;
data_inb = 16'h2;
#10;
address_ina = 202;
address_inb = 203;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 204;
address_inb = 205;
data_ina = 16'hffff;
data_inb = 16'hfffe;
#10;
address_ina = 206;
address_inb = 207;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 208;
address_inb = 209;
data_ina = 16'h0;
data_inb = 16'h3;
#10;
address_ina = 210;
address_inb = 211;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 212;
address_inb = 213;
data_ina = 16'hfffe;
data_inb = 16'h0;
#10;
address_ina = 214;
address_inb = 215;
data_ina = 16'h2;
data_inb = 16'h1;
#10;
address_ina = 216;
address_inb = 217;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 218;
address_inb = 219;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 220;
address_inb = 221;
data_ina = 16'h1;
data_inb = 16'h2;
#10;
address_ina = 222;
address_inb = 223;
data_ina = 16'h1;
data_inb = 16'h3;
#10;
address_ina = 224;
address_inb = 225;
data_ina = 16'h0;
data_inb = 16'hfffe;
#10;
address_ina = 226;
address_inb = 227;
data_ina = 16'hffff;
data_inb = 16'hfffe;
#10;
address_ina = 228;
address_inb = 229;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 230;
address_inb = 231;
data_ina = 16'h0;
data_inb = 16'h2;
#10;
address_ina = 232;
address_inb = 233;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 234;
address_inb = 235;
data_ina = 16'h0;
data_inb = 16'hfffe;
#10;
address_ina = 236;
address_inb = 237;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 238;
address_inb = 239;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 240;
address_inb = 241;
data_ina = 16'h2;
data_inb = 16'h1;
#10;
address_ina = 242;
address_inb = 243;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 244;
address_inb = 245;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 246;
address_inb = 247;
data_ina = 16'h1;
data_inb = 16'hfffd;
#10;
address_ina = 248;
address_inb = 249;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 250;
address_inb = 251;
data_ina = 16'h0;
data_inb = 16'hfffe;
#10;
address_ina = 252;
address_inb = 253;
data_ina = 16'h3;
data_inb = 16'hffff;
#10;
address_ina = 254;
address_inb = 255;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
        wait(init_done);
        #30
        we = 0;
        // Start processing
         
		  #38000

        start = 0;



//        wait (wr_req);
//		  wait (!wr_req);
//		   rd_req = 1;
		  wait(done);
		  #20000
rd_req = 1;
        #70 
		  start = 1;
		 #80 
wait(rd_empty)
rd_req = 0;

$display("Finished the NTT test Number %d",test_num);
////Begin test number #89//////////////
rst = 1;

//#1000
start = 1;
mode = 0; //NTT 0 // INTT 1

// Reset for a few clock cycles

#1000

rst = 0;
test_num = test_num + 1;
#1000
we = 1;
address_ina = 0;
address_inb = 1;
data_ina = 16'hfffe;
data_inb = 16'h0;
#10;
address_ina = 2;
address_inb = 3;
data_ina = 16'hffff;
data_inb = 16'hfffd;
#10;
address_ina = 4;
address_inb = 5;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 6;
address_inb = 7;
data_ina = 16'hfffe;
data_inb = 16'h1;
#10;
address_ina = 8;
address_inb = 9;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 10;
address_inb = 11;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 12;
address_inb = 13;
data_ina = 16'h3;
data_inb = 16'h1;
#10;
address_ina = 14;
address_inb = 15;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 16;
address_inb = 17;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 18;
address_inb = 19;
data_ina = 16'hffff;
data_inb = 16'h2;
#10;
address_ina = 20;
address_inb = 21;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 22;
address_inb = 23;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 24;
address_inb = 25;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 26;
address_inb = 27;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 28;
address_inb = 29;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 30;
address_inb = 31;
data_ina = 16'hfffe;
data_inb = 16'hffff;
#10;
address_ina = 32;
address_inb = 33;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 34;
address_inb = 35;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 36;
address_inb = 37;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 38;
address_inb = 39;
data_ina = 16'hfffe;
data_inb = 16'h1;
#10;
address_ina = 40;
address_inb = 41;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 42;
address_inb = 43;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 44;
address_inb = 45;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 46;
address_inb = 47;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 48;
address_inb = 49;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 50;
address_inb = 51;
data_ina = 16'h1;
data_inb = 16'hfffe;
#10;
address_ina = 52;
address_inb = 53;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 54;
address_inb = 55;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 56;
address_inb = 57;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 58;
address_inb = 59;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 60;
address_inb = 61;
data_ina = 16'hfffe;
data_inb = 16'h1;
#10;
address_ina = 62;
address_inb = 63;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 64;
address_inb = 65;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 66;
address_inb = 67;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 68;
address_inb = 69;
data_ina = 16'hffff;
data_inb = 16'hfffe;
#10;
address_ina = 70;
address_inb = 71;
data_ina = 16'h1;
data_inb = 16'hfffd;
#10;
address_ina = 72;
address_inb = 73;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 74;
address_inb = 75;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 76;
address_inb = 77;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 78;
address_inb = 79;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 80;
address_inb = 81;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 82;
address_inb = 83;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 84;
address_inb = 85;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 86;
address_inb = 87;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 88;
address_inb = 89;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 90;
address_inb = 91;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 92;
address_inb = 93;
data_ina = 16'h0;
data_inb = 16'hfffd;
#10;
address_ina = 94;
address_inb = 95;
data_ina = 16'h3;
data_inb = 16'h0;
#10;
address_ina = 96;
address_inb = 97;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 98;
address_inb = 99;
data_ina = 16'h1;
data_inb = 16'hfffe;
#10;
address_ina = 100;
address_inb = 101;
data_ina = 16'hfffd;
data_inb = 16'h0;
#10;
address_ina = 102;
address_inb = 103;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 104;
address_inb = 105;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 106;
address_inb = 107;
data_ina = 16'h2;
data_inb = 16'hffff;
#10;
address_ina = 108;
address_inb = 109;
data_ina = 16'hfffe;
data_inb = 16'hffff;
#10;
address_ina = 110;
address_inb = 111;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 112;
address_inb = 113;
data_ina = 16'hfffe;
data_inb = 16'hffff;
#10;
address_ina = 114;
address_inb = 115;
data_ina = 16'hfffd;
data_inb = 16'hffff;
#10;
address_ina = 116;
address_inb = 117;
data_ina = 16'hffff;
data_inb = 16'h3;
#10;
address_ina = 118;
address_inb = 119;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 120;
address_inb = 121;
data_ina = 16'h2;
data_inb = 16'hfffe;
#10;
address_ina = 122;
address_inb = 123;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 124;
address_inb = 125;
data_ina = 16'h2;
data_inb = 16'hffff;
#10;
address_ina = 126;
address_inb = 127;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 128;
address_inb = 129;
data_ina = 16'hfffd;
data_inb = 16'h2;
#10;
address_ina = 130;
address_inb = 131;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 132;
address_inb = 133;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 134;
address_inb = 135;
data_ina = 16'hfffe;
data_inb = 16'hffff;
#10;
address_ina = 136;
address_inb = 137;
data_ina = 16'h0;
data_inb = 16'h2;
#10;
address_ina = 138;
address_inb = 139;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 140;
address_inb = 141;
data_ina = 16'h2;
data_inb = 16'h1;
#10;
address_ina = 142;
address_inb = 143;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 144;
address_inb = 145;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 146;
address_inb = 147;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 148;
address_inb = 149;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 150;
address_inb = 151;
data_ina = 16'h1;
data_inb = 16'hfffe;
#10;
address_ina = 152;
address_inb = 153;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 154;
address_inb = 155;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 156;
address_inb = 157;
data_ina = 16'h2;
data_inb = 16'h0;
#10;
address_ina = 158;
address_inb = 159;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 160;
address_inb = 161;
data_ina = 16'hffff;
data_inb = 16'hfffe;
#10;
address_ina = 162;
address_inb = 163;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 164;
address_inb = 165;
data_ina = 16'h2;
data_inb = 16'h0;
#10;
address_ina = 166;
address_inb = 167;
data_ina = 16'h0;
data_inb = 16'hfffe;
#10;
address_ina = 168;
address_inb = 169;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 170;
address_inb = 171;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 172;
address_inb = 173;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 174;
address_inb = 175;
data_ina = 16'hffff;
data_inb = 16'hfffe;
#10;
address_ina = 176;
address_inb = 177;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 178;
address_inb = 179;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 180;
address_inb = 181;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 182;
address_inb = 183;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 184;
address_inb = 185;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 186;
address_inb = 187;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 188;
address_inb = 189;
data_ina = 16'h2;
data_inb = 16'h0;
#10;
address_ina = 190;
address_inb = 191;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 192;
address_inb = 193;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 194;
address_inb = 195;
data_ina = 16'h2;
data_inb = 16'h1;
#10;
address_ina = 196;
address_inb = 197;
data_ina = 16'h2;
data_inb = 16'h1;
#10;
address_ina = 198;
address_inb = 199;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 200;
address_inb = 201;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 202;
address_inb = 203;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 204;
address_inb = 205;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 206;
address_inb = 207;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 208;
address_inb = 209;
data_ina = 16'hffff;
data_inb = 16'hfffe;
#10;
address_ina = 210;
address_inb = 211;
data_ina = 16'h2;
data_inb = 16'h1;
#10;
address_ina = 212;
address_inb = 213;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 214;
address_inb = 215;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 216;
address_inb = 217;
data_ina = 16'h1;
data_inb = 16'h2;
#10;
address_ina = 218;
address_inb = 219;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 220;
address_inb = 221;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 222;
address_inb = 223;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 224;
address_inb = 225;
data_ina = 16'hffff;
data_inb = 16'hfffe;
#10;
address_ina = 226;
address_inb = 227;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 228;
address_inb = 229;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 230;
address_inb = 231;
data_ina = 16'hfffd;
data_inb = 16'hffff;
#10;
address_ina = 232;
address_inb = 233;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 234;
address_inb = 235;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 236;
address_inb = 237;
data_ina = 16'h1;
data_inb = 16'hfffe;
#10;
address_ina = 238;
address_inb = 239;
data_ina = 16'hfffe;
data_inb = 16'hffff;
#10;
address_ina = 240;
address_inb = 241;
data_ina = 16'hfffe;
data_inb = 16'hffff;
#10;
address_ina = 242;
address_inb = 243;
data_ina = 16'h1;
data_inb = 16'hfffe;
#10;
address_ina = 244;
address_inb = 245;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 246;
address_inb = 247;
data_ina = 16'hfffe;
data_inb = 16'h1;
#10;
address_ina = 248;
address_inb = 249;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 250;
address_inb = 251;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 252;
address_inb = 253;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 254;
address_inb = 255;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
        wait(init_done);
        #30
        we = 0;
        // Start processing
         
		  #38000

        start = 0;



//        wait (wr_req);
//		  wait (!wr_req);
//		   rd_req = 1;
		  wait(done);
		  #20000
rd_req = 1;
        #70 
		  start = 1;
		 #80 
wait(rd_empty)
rd_req = 0;

$display("Finished the NTT test Number %d",test_num);
////Begin test number #90//////////////
rst = 1;

//#1000
start = 1;
mode = 0; //NTT 0 // INTT 1

// Reset for a few clock cycles

#1000

rst = 0;
test_num = test_num + 1;
#1000
we = 1;
address_ina = 0;
address_inb = 1;
data_ina = 16'h2;
data_inb = 16'h1;
#10;
address_ina = 2;
address_inb = 3;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 4;
address_inb = 5;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 6;
address_inb = 7;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 8;
address_inb = 9;
data_ina = 16'hffff;
data_inb = 16'h2;
#10;
address_ina = 10;
address_inb = 11;
data_ina = 16'hffff;
data_inb = 16'h2;
#10;
address_ina = 12;
address_inb = 13;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 14;
address_inb = 15;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 16;
address_inb = 17;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 18;
address_inb = 19;
data_ina = 16'hfffe;
data_inb = 16'h0;
#10;
address_ina = 20;
address_inb = 21;
data_ina = 16'hffff;
data_inb = 16'hfffe;
#10;
address_ina = 22;
address_inb = 23;
data_ina = 16'h3;
data_inb = 16'h0;
#10;
address_ina = 24;
address_inb = 25;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 26;
address_inb = 27;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 28;
address_inb = 29;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 30;
address_inb = 31;
data_ina = 16'hffff;
data_inb = 16'hfffe;
#10;
address_ina = 32;
address_inb = 33;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 34;
address_inb = 35;
data_ina = 16'hfffe;
data_inb = 16'hffff;
#10;
address_ina = 36;
address_inb = 37;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 38;
address_inb = 39;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 40;
address_inb = 41;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 42;
address_inb = 43;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 44;
address_inb = 45;
data_ina = 16'hffff;
data_inb = 16'hfffe;
#10;
address_ina = 46;
address_inb = 47;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 48;
address_inb = 49;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 50;
address_inb = 51;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 52;
address_inb = 53;
data_ina = 16'h2;
data_inb = 16'hfffe;
#10;
address_ina = 54;
address_inb = 55;
data_ina = 16'h0;
data_inb = 16'hfffe;
#10;
address_ina = 56;
address_inb = 57;
data_ina = 16'hfffe;
data_inb = 16'h0;
#10;
address_ina = 58;
address_inb = 59;
data_ina = 16'h1;
data_inb = 16'h2;
#10;
address_ina = 60;
address_inb = 61;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 62;
address_inb = 63;
data_ina = 16'hffff;
data_inb = 16'h2;
#10;
address_ina = 64;
address_inb = 65;
data_ina = 16'hfffe;
data_inb = 16'h0;
#10;
address_ina = 66;
address_inb = 67;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 68;
address_inb = 69;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 70;
address_inb = 71;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 72;
address_inb = 73;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 74;
address_inb = 75;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 76;
address_inb = 77;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 78;
address_inb = 79;
data_ina = 16'h1;
data_inb = 16'h2;
#10;
address_ina = 80;
address_inb = 81;
data_ina = 16'h2;
data_inb = 16'h3;
#10;
address_ina = 82;
address_inb = 83;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 84;
address_inb = 85;
data_ina = 16'hfffe;
data_inb = 16'hffff;
#10;
address_ina = 86;
address_inb = 87;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 88;
address_inb = 89;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 90;
address_inb = 91;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 92;
address_inb = 93;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 94;
address_inb = 95;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 96;
address_inb = 97;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 98;
address_inb = 99;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 100;
address_inb = 101;
data_ina = 16'h0;
data_inb = 16'h3;
#10;
address_ina = 102;
address_inb = 103;
data_ina = 16'h2;
data_inb = 16'h0;
#10;
address_ina = 104;
address_inb = 105;
data_ina = 16'hfffe;
data_inb = 16'h1;
#10;
address_ina = 106;
address_inb = 107;
data_ina = 16'hfffe;
data_inb = 16'hffff;
#10;
address_ina = 108;
address_inb = 109;
data_ina = 16'hfffe;
data_inb = 16'h0;
#10;
address_ina = 110;
address_inb = 111;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 112;
address_inb = 113;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 114;
address_inb = 115;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 116;
address_inb = 117;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 118;
address_inb = 119;
data_ina = 16'hfffd;
data_inb = 16'hfffe;
#10;
address_ina = 120;
address_inb = 121;
data_ina = 16'h1;
data_inb = 16'hfffe;
#10;
address_ina = 122;
address_inb = 123;
data_ina = 16'h1;
data_inb = 16'hfffe;
#10;
address_ina = 124;
address_inb = 125;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 126;
address_inb = 127;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 128;
address_inb = 129;
data_ina = 16'h1;
data_inb = 16'h3;
#10;
address_ina = 130;
address_inb = 131;
data_ina = 16'h0;
data_inb = 16'h2;
#10;
address_ina = 132;
address_inb = 133;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 134;
address_inb = 135;
data_ina = 16'h2;
data_inb = 16'h0;
#10;
address_ina = 136;
address_inb = 137;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 138;
address_inb = 139;
data_ina = 16'h0;
data_inb = 16'h2;
#10;
address_ina = 140;
address_inb = 141;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 142;
address_inb = 143;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 144;
address_inb = 145;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 146;
address_inb = 147;
data_ina = 16'hfffe;
data_inb = 16'h1;
#10;
address_ina = 148;
address_inb = 149;
data_ina = 16'hfffd;
data_inb = 16'h1;
#10;
address_ina = 150;
address_inb = 151;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 152;
address_inb = 153;
data_ina = 16'h2;
data_inb = 16'h2;
#10;
address_ina = 154;
address_inb = 155;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 156;
address_inb = 157;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 158;
address_inb = 159;
data_ina = 16'h2;
data_inb = 16'h3;
#10;
address_ina = 160;
address_inb = 161;
data_ina = 16'h2;
data_inb = 16'hffff;
#10;
address_ina = 162;
address_inb = 163;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 164;
address_inb = 165;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 166;
address_inb = 167;
data_ina = 16'hffff;
data_inb = 16'h3;
#10;
address_ina = 168;
address_inb = 169;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 170;
address_inb = 171;
data_ina = 16'h2;
data_inb = 16'hfffe;
#10;
address_ina = 172;
address_inb = 173;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 174;
address_inb = 175;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 176;
address_inb = 177;
data_ina = 16'h1;
data_inb = 16'h2;
#10;
address_ina = 178;
address_inb = 179;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 180;
address_inb = 181;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 182;
address_inb = 183;
data_ina = 16'h2;
data_inb = 16'hffff;
#10;
address_ina = 184;
address_inb = 185;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 186;
address_inb = 187;
data_ina = 16'hffff;
data_inb = 16'h2;
#10;
address_ina = 188;
address_inb = 189;
data_ina = 16'h3;
data_inb = 16'hffff;
#10;
address_ina = 190;
address_inb = 191;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 192;
address_inb = 193;
data_ina = 16'h0;
data_inb = 16'hfffe;
#10;
address_ina = 194;
address_inb = 195;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 196;
address_inb = 197;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 198;
address_inb = 199;
data_ina = 16'hfffe;
data_inb = 16'h0;
#10;
address_ina = 200;
address_inb = 201;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 202;
address_inb = 203;
data_ina = 16'h3;
data_inb = 16'h0;
#10;
address_ina = 204;
address_inb = 205;
data_ina = 16'h3;
data_inb = 16'h1;
#10;
address_ina = 206;
address_inb = 207;
data_ina = 16'h0;
data_inb = 16'hfffe;
#10;
address_ina = 208;
address_inb = 209;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 210;
address_inb = 211;
data_ina = 16'hfffe;
data_inb = 16'h0;
#10;
address_ina = 212;
address_inb = 213;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 214;
address_inb = 215;
data_ina = 16'h0;
data_inb = 16'h3;
#10;
address_ina = 216;
address_inb = 217;
data_ina = 16'hffff;
data_inb = 16'hfffe;
#10;
address_ina = 218;
address_inb = 219;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 220;
address_inb = 221;
data_ina = 16'h2;
data_inb = 16'h0;
#10;
address_ina = 222;
address_inb = 223;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 224;
address_inb = 225;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 226;
address_inb = 227;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 228;
address_inb = 229;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 230;
address_inb = 231;
data_ina = 16'hfffe;
data_inb = 16'h0;
#10;
address_ina = 232;
address_inb = 233;
data_ina = 16'hfffe;
data_inb = 16'h2;
#10;
address_ina = 234;
address_inb = 235;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 236;
address_inb = 237;
data_ina = 16'h0;
data_inb = 16'h2;
#10;
address_ina = 238;
address_inb = 239;
data_ina = 16'hfffd;
data_inb = 16'hfffe;
#10;
address_ina = 240;
address_inb = 241;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 242;
address_inb = 243;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 244;
address_inb = 245;
data_ina = 16'hfffe;
data_inb = 16'h0;
#10;
address_ina = 246;
address_inb = 247;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 248;
address_inb = 249;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 250;
address_inb = 251;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 252;
address_inb = 253;
data_ina = 16'hfffe;
data_inb = 16'h1;
#10;
address_ina = 254;
address_inb = 255;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
        wait(init_done);
        #30
        we = 0;
        // Start processing
         
		  #38000

        start = 0;



//        wait (wr_req);
//		  wait (!wr_req);
//		   rd_req = 1;
		  wait(done);
		  #20000
rd_req = 1;
        #70 
		  start = 1;
		 #80 
wait(rd_empty)
rd_req = 0;

$display("Finished the NTT test Number %d",test_num);
////Begin test number #91//////////////
rst = 1;

//#1000
start = 1;
mode = 1; //NTT 0 // INTT 1

// Reset for a few clock cycles

#1000

rst = 0;
test_num = test_num + 1;
#1000
we = 1;
address_ina = 0;
address_inb = 1;
data_ina = 16'h37f;
data_inb = 16'h5c3;
#10;
address_ina = 2;
address_inb = 3;
data_ina = 16'h313;
data_inb = 16'h233;
#10;
address_ina = 4;
address_inb = 5;
data_ina = 16'hf9d9;
data_inb = 16'h201;
#10;
address_ina = 6;
address_inb = 7;
data_ina = 16'h49b;
data_inb = 16'h9c;
#10;
address_ina = 8;
address_inb = 9;
data_ina = 16'h35b;
data_inb = 16'hf9cb;
#10;
address_ina = 10;
address_inb = 11;
data_ina = 16'hf98e;
data_inb = 16'h638;
#10;
address_ina = 12;
address_inb = 13;
data_ina = 16'h2c7;
data_inb = 16'h3a1;
#10;
address_ina = 14;
address_inb = 15;
data_ina = 16'h47c;
data_inb = 16'hfde5;
#10;
address_ina = 16;
address_inb = 17;
data_ina = 16'hff6f;
data_inb = 16'h3d4;
#10;
address_ina = 18;
address_inb = 19;
data_ina = 16'h299;
data_inb = 16'hff45;
#10;
address_ina = 20;
address_inb = 21;
data_ina = 16'hfd26;
data_inb = 16'hfb12;
#10;
address_ina = 22;
address_inb = 23;
data_ina = 16'hfb51;
data_inb = 16'hfe5d;
#10;
address_ina = 24;
address_inb = 25;
data_ina = 16'hfbf7;
data_inb = 16'h383;
#10;
address_ina = 26;
address_inb = 27;
data_ina = 16'hfb14;
data_inb = 16'h47;
#10;
address_ina = 28;
address_inb = 29;
data_ina = 16'h98;
data_inb = 16'hff1a;
#10;
address_ina = 30;
address_inb = 31;
data_ina = 16'h1b2;
data_inb = 16'h202;
#10;
address_ina = 32;
address_inb = 33;
data_ina = 16'hfb27;
data_inb = 16'h5c8;
#10;
address_ina = 34;
address_inb = 35;
data_ina = 16'h454;
data_inb = 16'h4c8;
#10;
address_ina = 36;
address_inb = 37;
data_ina = 16'hffea;
data_inb = 16'h2f0;
#10;
address_ina = 38;
address_inb = 39;
data_ina = 16'h3d1;
data_inb = 16'h3c9;
#10;
address_ina = 40;
address_inb = 41;
data_ina = 16'h51c;
data_inb = 16'hfb5b;
#10;
address_ina = 42;
address_inb = 43;
data_ina = 16'hfd3e;
data_inb = 16'hfa35;
#10;
address_ina = 44;
address_inb = 45;
data_ina = 16'h492;
data_inb = 16'h18f;
#10;
address_ina = 46;
address_inb = 47;
data_ina = 16'hfb19;
data_inb = 16'h259;
#10;
address_ina = 48;
address_inb = 49;
data_ina = 16'hfd2a;
data_inb = 16'h5be;
#10;
address_ina = 50;
address_inb = 51;
data_ina = 16'hfc9f;
data_inb = 16'hff19;
#10;
address_ina = 52;
address_inb = 53;
data_ina = 16'h26b;
data_inb = 16'hfedf;
#10;
address_ina = 54;
address_inb = 55;
data_ina = 16'hfa74;
data_inb = 16'hfcf5;
#10;
address_ina = 56;
address_inb = 57;
data_ina = 16'hfe2a;
data_inb = 16'h5ab;
#10;
address_ina = 58;
address_inb = 59;
data_ina = 16'h21f;
data_inb = 16'h413;
#10;
address_ina = 60;
address_inb = 61;
data_ina = 16'hfa24;
data_inb = 16'h67b;
#10;
address_ina = 62;
address_inb = 63;
data_ina = 16'h13b;
data_inb = 16'h620;
#10;
address_ina = 64;
address_inb = 65;
data_ina = 16'h6c;
data_inb = 16'hfd4e;
#10;
address_ina = 66;
address_inb = 67;
data_ina = 16'h262;
data_inb = 16'h56a;
#10;
address_ina = 68;
address_inb = 69;
data_ina = 16'hfc16;
data_inb = 16'hfda0;
#10;
address_ina = 70;
address_inb = 71;
data_ina = 16'h81;
data_inb = 16'h1bd;
#10;
address_ina = 72;
address_inb = 73;
data_ina = 16'h28a;
data_inb = 16'h31c;
#10;
address_ina = 74;
address_inb = 75;
data_ina = 16'hfde2;
data_inb = 16'hf9f0;
#10;
address_ina = 76;
address_inb = 77;
data_ina = 16'h46d;
data_inb = 16'hfd1c;
#10;
address_ina = 78;
address_inb = 79;
data_ina = 16'hff92;
data_inb = 16'hfa31;
#10;
address_ina = 80;
address_inb = 81;
data_ina = 16'h3f0;
data_inb = 16'hfd75;
#10;
address_ina = 82;
address_inb = 83;
data_ina = 16'h3;
data_inb = 16'h4c8;
#10;
address_ina = 84;
address_inb = 85;
data_ina = 16'hff72;
data_inb = 16'hfb9a;
#10;
address_ina = 86;
address_inb = 87;
data_ina = 16'hfe33;
data_inb = 16'h674;
#10;
address_ina = 88;
address_inb = 89;
data_ina = 16'hfd41;
data_inb = 16'hfdb8;
#10;
address_ina = 90;
address_inb = 91;
data_ina = 16'h2d2;
data_inb = 16'h4ed;
#10;
address_ina = 92;
address_inb = 93;
data_ina = 16'hfa49;
data_inb = 16'h625;
#10;
address_ina = 94;
address_inb = 95;
data_ina = 16'h358;
data_inb = 16'hfc86;
#10;
address_ina = 96;
address_inb = 97;
data_ina = 16'h3b;
data_inb = 16'h4ba;
#10;
address_ina = 98;
address_inb = 99;
data_ina = 16'h5e1;
data_inb = 16'h27c;
#10;
address_ina = 100;
address_inb = 101;
data_ina = 16'hfcc5;
data_inb = 16'h47c;
#10;
address_ina = 102;
address_inb = 103;
data_ina = 16'hfd11;
data_inb = 16'h5a1;
#10;
address_ina = 104;
address_inb = 105;
data_ina = 16'hfebd;
data_inb = 16'h3d6;
#10;
address_ina = 106;
address_inb = 107;
data_ina = 16'hffbe;
data_inb = 16'hf9e6;
#10;
address_ina = 108;
address_inb = 109;
data_ina = 16'h2ad;
data_inb = 16'h1df;
#10;
address_ina = 110;
address_inb = 111;
data_ina = 16'h642;
data_inb = 16'hf9ba;
#10;
address_ina = 112;
address_inb = 113;
data_ina = 16'hf9eb;
data_inb = 16'h235;
#10;
address_ina = 114;
address_inb = 115;
data_ina = 16'h223;
data_inb = 16'hfe7e;
#10;
address_ina = 116;
address_inb = 117;
data_ina = 16'h20b;
data_inb = 16'hfc43;
#10;
address_ina = 118;
address_inb = 119;
data_ina = 16'h633;
data_inb = 16'h48c;
#10;
address_ina = 120;
address_inb = 121;
data_ina = 16'hfd47;
data_inb = 16'h19d;
#10;
address_ina = 122;
address_inb = 123;
data_ina = 16'h515;
data_inb = 16'hc8;
#10;
address_ina = 124;
address_inb = 125;
data_ina = 16'hfa09;
data_inb = 16'h78;
#10;
address_ina = 126;
address_inb = 127;
data_ina = 16'h9;
data_inb = 16'h177;
#10;
address_ina = 128;
address_inb = 129;
data_ina = 16'h41b;
data_inb = 16'h11b;
#10;
address_ina = 130;
address_inb = 131;
data_ina = 16'hfb8d;
data_inb = 16'hfe3d;
#10;
address_ina = 132;
address_inb = 133;
data_ina = 16'hfbc5;
data_inb = 16'h23;
#10;
address_ina = 134;
address_inb = 135;
data_ina = 16'hfd81;
data_inb = 16'h12;
#10;
address_ina = 136;
address_inb = 137;
data_ina = 16'hfc86;
data_inb = 16'hfaa2;
#10;
address_ina = 138;
address_inb = 139;
data_ina = 16'h39f;
data_inb = 16'h16f;
#10;
address_ina = 140;
address_inb = 141;
data_ina = 16'hfc19;
data_inb = 16'hf9b9;
#10;
address_ina = 142;
address_inb = 143;
data_ina = 16'h27;
data_inb = 16'he3;
#10;
address_ina = 144;
address_inb = 145;
data_ina = 16'h3f1;
data_inb = 16'h72;
#10;
address_ina = 146;
address_inb = 147;
data_ina = 16'hfe51;
data_inb = 16'hfeb0;
#10;
address_ina = 148;
address_inb = 149;
data_ina = 16'h604;
data_inb = 16'h317;
#10;
address_ina = 150;
address_inb = 151;
data_ina = 16'hfa15;
data_inb = 16'hfb77;
#10;
address_ina = 152;
address_inb = 153;
data_ina = 16'h3bf;
data_inb = 16'h21f;
#10;
address_ina = 154;
address_inb = 155;
data_ina = 16'h3a4;
data_inb = 16'hfd53;
#10;
address_ina = 156;
address_inb = 157;
data_ina = 16'h4c4;
data_inb = 16'hfd7b;
#10;
address_ina = 158;
address_inb = 159;
data_ina = 16'h17a;
data_inb = 16'hf7;
#10;
address_ina = 160;
address_inb = 161;
data_ina = 16'h313;
data_inb = 16'h2a5;
#10;
address_ina = 162;
address_inb = 163;
data_ina = 16'hfcc2;
data_inb = 16'hfa44;
#10;
address_ina = 164;
address_inb = 165;
data_ina = 16'h4c3;
data_inb = 16'h4c0;
#10;
address_ina = 166;
address_inb = 167;
data_ina = 16'hfdc8;
data_inb = 16'hfe5d;
#10;
address_ina = 168;
address_inb = 169;
data_ina = 16'hf9ce;
data_inb = 16'hf9e4;
#10;
address_ina = 170;
address_inb = 171;
data_ina = 16'h4;
data_inb = 16'hfbd4;
#10;
address_ina = 172;
address_inb = 173;
data_ina = 16'h443;
data_inb = 16'h49d;
#10;
address_ina = 174;
address_inb = 175;
data_ina = 16'hfd64;
data_inb = 16'hfeda;
#10;
address_ina = 176;
address_inb = 177;
data_ina = 16'hf9c8;
data_inb = 16'hff4f;
#10;
address_ina = 178;
address_inb = 179;
data_ina = 16'hfeec;
data_inb = 16'hff92;
#10;
address_ina = 180;
address_inb = 181;
data_ina = 16'hfde3;
data_inb = 16'hfe9e;
#10;
address_ina = 182;
address_inb = 183;
data_ina = 16'haa;
data_inb = 16'hfafa;
#10;
address_ina = 184;
address_inb = 185;
data_ina = 16'hf9aa;
data_inb = 16'h623;
#10;
address_ina = 186;
address_inb = 187;
data_ina = 16'h14a;
data_inb = 16'hfd50;
#10;
address_ina = 188;
address_inb = 189;
data_ina = 16'h53a;
data_inb = 16'h24b;
#10;
address_ina = 190;
address_inb = 191;
data_ina = 16'h33f;
data_inb = 16'h280;
#10;
address_ina = 192;
address_inb = 193;
data_ina = 16'h187;
data_inb = 16'h35c;
#10;
address_ina = 194;
address_inb = 195;
data_ina = 16'hfd97;
data_inb = 16'h3b6;
#10;
address_ina = 196;
address_inb = 197;
data_ina = 16'hfa4f;
data_inb = 16'h240;
#10;
address_ina = 198;
address_inb = 199;
data_ina = 16'hfd2c;
data_inb = 16'hff50;
#10;
address_ina = 200;
address_inb = 201;
data_ina = 16'h2ad;
data_inb = 16'h5d4;
#10;
address_ina = 202;
address_inb = 203;
data_ina = 16'h60c;
data_inb = 16'hfda3;
#10;
address_ina = 204;
address_inb = 205;
data_ina = 16'h144;
data_inb = 16'h2fc;
#10;
address_ina = 206;
address_inb = 207;
data_ina = 16'h197;
data_inb = 16'h370;
#10;
address_ina = 208;
address_inb = 209;
data_ina = 16'h590;
data_inb = 16'h44a;
#10;
address_ina = 210;
address_inb = 211;
data_ina = 16'hfffd;
data_inb = 16'h83;
#10;
address_ina = 212;
address_inb = 213;
data_ina = 16'hfff8;
data_inb = 16'h2c2;
#10;
address_ina = 214;
address_inb = 215;
data_ina = 16'h8f;
data_inb = 16'h228;
#10;
address_ina = 216;
address_inb = 217;
data_ina = 16'h224;
data_inb = 16'hfcd5;
#10;
address_ina = 218;
address_inb = 219;
data_ina = 16'h586;
data_inb = 16'h123;
#10;
address_ina = 220;
address_inb = 221;
data_ina = 16'hf9ce;
data_inb = 16'h268;
#10;
address_ina = 222;
address_inb = 223;
data_ina = 16'h516;
data_inb = 16'h558;
#10;
address_ina = 224;
address_inb = 225;
data_ina = 16'h1a1;
data_inb = 16'hfa5d;
#10;
address_ina = 226;
address_inb = 227;
data_ina = 16'hfe7d;
data_inb = 16'hfce2;
#10;
address_ina = 228;
address_inb = 229;
data_ina = 16'hfeaa;
data_inb = 16'hfb2b;
#10;
address_ina = 230;
address_inb = 231;
data_ina = 16'hfdad;
data_inb = 16'h22;
#10;
address_ina = 232;
address_inb = 233;
data_ina = 16'hd3;
data_inb = 16'hff95;
#10;
address_ina = 234;
address_inb = 235;
data_ina = 16'h437;
data_inb = 16'hfbf8;
#10;
address_ina = 236;
address_inb = 237;
data_ina = 16'h51f;
data_inb = 16'hfbda;
#10;
address_ina = 238;
address_inb = 239;
data_ina = 16'hfc4d;
data_inb = 16'h4cf;
#10;
address_ina = 240;
address_inb = 241;
data_ina = 16'hfcbc;
data_inb = 16'hfd8f;
#10;
address_ina = 242;
address_inb = 243;
data_ina = 16'h41c;
data_inb = 16'hfe2f;
#10;
address_ina = 244;
address_inb = 245;
data_ina = 16'hfa24;
data_inb = 16'hfe58;
#10;
address_ina = 246;
address_inb = 247;
data_ina = 16'hfe6a;
data_inb = 16'hfc2c;
#10;
address_ina = 248;
address_inb = 249;
data_ina = 16'h469;
data_inb = 16'hfd84;
#10;
address_ina = 250;
address_inb = 251;
data_ina = 16'hf9c6;
data_inb = 16'hfc46;
#10;
address_ina = 252;
address_inb = 253;
data_ina = 16'hfc73;
data_inb = 16'hfdce;
#10;
address_ina = 254;
address_inb = 255;
data_ina = 16'h3d5;
data_inb = 16'hfc99;
#10;
        wait(init_done);
        #30
        we = 0;
        // Start processing
         
		  #38000

        start = 0;



//        wait (wr_req);
//		  wait (!wr_req);
//		   rd_req = 1;
		  wait(done);
		  #20000
rd_req = 1;
        #70 
		  start = 1;
		 #80 
wait(rd_empty)
rd_req = 0;

$display("Finished the NTT test Number %d",test_num);
////Begin test number #92//////////////
rst = 1;

//#1000
start = 1;
mode = 1; //NTT 0 // INTT 1

// Reset for a few clock cycles

#1000

rst = 0;
test_num = test_num + 1;
#1000
we = 1;
address_ina = 0;
address_inb = 1;
data_ina = 16'h18f;
data_inb = 16'h3c3;
#10;
address_ina = 2;
address_inb = 3;
data_ina = 16'hfbda;
data_inb = 16'hfde0;
#10;
address_ina = 4;
address_inb = 5;
data_ina = 16'h3a3;
data_inb = 16'hfc7e;
#10;
address_ina = 6;
address_inb = 7;
data_ina = 16'h557;
data_inb = 16'hfc18;
#10;
address_ina = 8;
address_inb = 9;
data_ina = 16'h590;
data_inb = 16'hfa2c;
#10;
address_ina = 10;
address_inb = 11;
data_ina = 16'h5a1;
data_inb = 16'hf9a4;
#10;
address_ina = 12;
address_inb = 13;
data_ina = 16'h8;
data_inb = 16'h16e;
#10;
address_ina = 14;
address_inb = 15;
data_ina = 16'hff62;
data_inb = 16'hfcc1;
#10;
address_ina = 16;
address_inb = 17;
data_ina = 16'h2de;
data_inb = 16'hff88;
#10;
address_ina = 18;
address_inb = 19;
data_ina = 16'h163;
data_inb = 16'hfb1e;
#10;
address_ina = 20;
address_inb = 21;
data_ina = 16'h152;
data_inb = 16'hfd25;
#10;
address_ina = 22;
address_inb = 23;
data_ina = 16'hfdc5;
data_inb = 16'h5b0;
#10;
address_ina = 24;
address_inb = 25;
data_ina = 16'h3b5;
data_inb = 16'h66f;
#10;
address_ina = 26;
address_inb = 27;
data_ina = 16'h5e2;
data_inb = 16'hff61;
#10;
address_ina = 28;
address_inb = 29;
data_ina = 16'h36c;
data_inb = 16'h37b;
#10;
address_ina = 30;
address_inb = 31;
data_ina = 16'hfaba;
data_inb = 16'hfb53;
#10;
address_ina = 32;
address_inb = 33;
data_ina = 16'hfec5;
data_inb = 16'hff54;
#10;
address_ina = 34;
address_inb = 35;
data_ina = 16'hfa55;
data_inb = 16'h3e;
#10;
address_ina = 36;
address_inb = 37;
data_ina = 16'h5ce;
data_inb = 16'hffb6;
#10;
address_ina = 38;
address_inb = 39;
data_ina = 16'hff17;
data_inb = 16'hf9e2;
#10;
address_ina = 40;
address_inb = 41;
data_ina = 16'hce;
data_inb = 16'hf9b0;
#10;
address_ina = 42;
address_inb = 43;
data_ina = 16'h1e0;
data_inb = 16'h639;
#10;
address_ina = 44;
address_inb = 45;
data_ina = 16'h4f5;
data_inb = 16'h9f;
#10;
address_ina = 46;
address_inb = 47;
data_ina = 16'h46a;
data_inb = 16'hf99d;
#10;
address_ina = 48;
address_inb = 49;
data_ina = 16'h3e6;
data_inb = 16'hff9d;
#10;
address_ina = 50;
address_inb = 51;
data_ina = 16'hfa67;
data_inb = 16'h660;
#10;
address_ina = 52;
address_inb = 53;
data_ina = 16'hfcac;
data_inb = 16'h45f;
#10;
address_ina = 54;
address_inb = 55;
data_ina = 16'h65;
data_inb = 16'h52c;
#10;
address_ina = 56;
address_inb = 57;
data_ina = 16'hfc14;
data_inb = 16'h452;
#10;
address_ina = 58;
address_inb = 59;
data_ina = 16'hffd2;
data_inb = 16'hfc5d;
#10;
address_ina = 60;
address_inb = 61;
data_ina = 16'hfc4a;
data_inb = 16'hfd29;
#10;
address_ina = 62;
address_inb = 63;
data_ina = 16'h234;
data_inb = 16'hfddb;
#10;
address_ina = 64;
address_inb = 65;
data_ina = 16'hfe41;
data_inb = 16'h269;
#10;
address_ina = 66;
address_inb = 67;
data_ina = 16'hfb24;
data_inb = 16'hfd60;
#10;
address_ina = 68;
address_inb = 69;
data_ina = 16'hf5;
data_inb = 16'h406;
#10;
address_ina = 70;
address_inb = 71;
data_ina = 16'h11b;
data_inb = 16'h504;
#10;
address_ina = 72;
address_inb = 73;
data_ina = 16'hfe7c;
data_inb = 16'hfbae;
#10;
address_ina = 74;
address_inb = 75;
data_ina = 16'hff64;
data_inb = 16'hfd7c;
#10;
address_ina = 76;
address_inb = 77;
data_ina = 16'h63e;
data_inb = 16'hfad8;
#10;
address_ina = 78;
address_inb = 79;
data_ina = 16'h3c5;
data_inb = 16'h19d;
#10;
address_ina = 80;
address_inb = 81;
data_ina = 16'hfb86;
data_inb = 16'h66a;
#10;
address_ina = 82;
address_inb = 83;
data_ina = 16'hfb29;
data_inb = 16'hfd4a;
#10;
address_ina = 84;
address_inb = 85;
data_ina = 16'hfcd8;
data_inb = 16'hfb78;
#10;
address_ina = 86;
address_inb = 87;
data_ina = 16'h2fe;
data_inb = 16'h4c4;
#10;
address_ina = 88;
address_inb = 89;
data_ina = 16'hfa5f;
data_inb = 16'h5ce;
#10;
address_ina = 90;
address_inb = 91;
data_ina = 16'h1ee;
data_inb = 16'hfbd7;
#10;
address_ina = 92;
address_inb = 93;
data_ina = 16'hfaec;
data_inb = 16'h2c4;
#10;
address_ina = 94;
address_inb = 95;
data_ina = 16'hfde2;
data_inb = 16'h42d;
#10;
address_ina = 96;
address_inb = 97;
data_ina = 16'hfef5;
data_inb = 16'h58f;
#10;
address_ina = 98;
address_inb = 99;
data_ina = 16'hf9cc;
data_inb = 16'hff46;
#10;
address_ina = 100;
address_inb = 101;
data_ina = 16'h496;
data_inb = 16'h45c;
#10;
address_ina = 102;
address_inb = 103;
data_ina = 16'hfe22;
data_inb = 16'h610;
#10;
address_ina = 104;
address_inb = 105;
data_ina = 16'h34e;
data_inb = 16'h4c1;
#10;
address_ina = 106;
address_inb = 107;
data_ina = 16'hf982;
data_inb = 16'hfff1;
#10;
address_ina = 108;
address_inb = 109;
data_ina = 16'hfef6;
data_inb = 16'hfcc7;
#10;
address_ina = 110;
address_inb = 111;
data_ina = 16'h173;
data_inb = 16'hfc7a;
#10;
address_ina = 112;
address_inb = 113;
data_ina = 16'ha1;
data_inb = 16'hff79;
#10;
address_ina = 114;
address_inb = 115;
data_ina = 16'h3dd;
data_inb = 16'h54a;
#10;
address_ina = 116;
address_inb = 117;
data_ina = 16'hfa68;
data_inb = 16'h4c3;
#10;
address_ina = 118;
address_inb = 119;
data_ina = 16'hfa7e;
data_inb = 16'h505;
#10;
address_ina = 120;
address_inb = 121;
data_ina = 16'h55a;
data_inb = 16'h2c7;
#10;
address_ina = 122;
address_inb = 123;
data_ina = 16'hfe00;
data_inb = 16'h1cd;
#10;
address_ina = 124;
address_inb = 125;
data_ina = 16'hff31;
data_inb = 16'hfe8f;
#10;
address_ina = 126;
address_inb = 127;
data_ina = 16'hfc3c;
data_inb = 16'hfbd1;
#10;
address_ina = 128;
address_inb = 129;
data_ina = 16'h54f;
data_inb = 16'h38;
#10;
address_ina = 130;
address_inb = 131;
data_ina = 16'h2f3;
data_inb = 16'h48d;
#10;
address_ina = 132;
address_inb = 133;
data_ina = 16'hffde;
data_inb = 16'h414;
#10;
address_ina = 134;
address_inb = 135;
data_ina = 16'h205;
data_inb = 16'hf9ed;
#10;
address_ina = 136;
address_inb = 137;
data_ina = 16'hfce0;
data_inb = 16'h653;
#10;
address_ina = 138;
address_inb = 139;
data_ina = 16'h26e;
data_inb = 16'hfcf1;
#10;
address_ina = 140;
address_inb = 141;
data_ina = 16'h192;
data_inb = 16'hfa43;
#10;
address_ina = 142;
address_inb = 143;
data_ina = 16'hfefc;
data_inb = 16'h89;
#10;
address_ina = 144;
address_inb = 145;
data_ina = 16'h486;
data_inb = 16'hfa5a;
#10;
address_ina = 146;
address_inb = 147;
data_ina = 16'h2ca;
data_inb = 16'h514;
#10;
address_ina = 148;
address_inb = 149;
data_ina = 16'h8c;
data_inb = 16'hffc8;
#10;
address_ina = 150;
address_inb = 151;
data_ina = 16'h2c7;
data_inb = 16'hfa6d;
#10;
address_ina = 152;
address_inb = 153;
data_ina = 16'hfc2e;
data_inb = 16'hfc0f;
#10;
address_ina = 154;
address_inb = 155;
data_ina = 16'hfd63;
data_inb = 16'h4ae;
#10;
address_ina = 156;
address_inb = 157;
data_ina = 16'hfbc4;
data_inb = 16'hfa08;
#10;
address_ina = 158;
address_inb = 159;
data_ina = 16'h350;
data_inb = 16'hfe10;
#10;
address_ina = 160;
address_inb = 161;
data_ina = 16'h471;
data_inb = 16'hfbf8;
#10;
address_ina = 162;
address_inb = 163;
data_ina = 16'hfa9f;
data_inb = 16'h353;
#10;
address_ina = 164;
address_inb = 165;
data_ina = 16'h342;
data_inb = 16'hfaba;
#10;
address_ina = 166;
address_inb = 167;
data_ina = 16'h4ad;
data_inb = 16'h26a;
#10;
address_ina = 168;
address_inb = 169;
data_ina = 16'hfc1b;
data_inb = 16'h213;
#10;
address_ina = 170;
address_inb = 171;
data_ina = 16'h1c0;
data_inb = 16'h271;
#10;
address_ina = 172;
address_inb = 173;
data_ina = 16'hf7;
data_inb = 16'hfec8;
#10;
address_ina = 174;
address_inb = 175;
data_ina = 16'h2db;
data_inb = 16'hf2;
#10;
address_ina = 176;
address_inb = 177;
data_ina = 16'hfe44;
data_inb = 16'hfa80;
#10;
address_ina = 178;
address_inb = 179;
data_ina = 16'h130;
data_inb = 16'h34f;
#10;
address_ina = 180;
address_inb = 181;
data_ina = 16'h470;
data_inb = 16'hfee0;
#10;
address_ina = 182;
address_inb = 183;
data_ina = 16'hfbc4;
data_inb = 16'h665;
#10;
address_ina = 184;
address_inb = 185;
data_ina = 16'h24d;
data_inb = 16'h170;
#10;
address_ina = 186;
address_inb = 187;
data_ina = 16'h4db;
data_inb = 16'hffc8;
#10;
address_ina = 188;
address_inb = 189;
data_ina = 16'h2ae;
data_inb = 16'hfbd0;
#10;
address_ina = 190;
address_inb = 191;
data_ina = 16'hfa2d;
data_inb = 16'hf98e;
#10;
address_ina = 192;
address_inb = 193;
data_ina = 16'h577;
data_inb = 16'h55e;
#10;
address_ina = 194;
address_inb = 195;
data_ina = 16'hfeac;
data_inb = 16'h60e;
#10;
address_ina = 196;
address_inb = 197;
data_ina = 16'hffe9;
data_inb = 16'h415;
#10;
address_ina = 198;
address_inb = 199;
data_ina = 16'hfb51;
data_inb = 16'h1a6;
#10;
address_ina = 200;
address_inb = 201;
data_ina = 16'hff96;
data_inb = 16'hfa73;
#10;
address_ina = 202;
address_inb = 203;
data_ina = 16'hfd2d;
data_inb = 16'hfad5;
#10;
address_ina = 204;
address_inb = 205;
data_ina = 16'hf9d8;
data_inb = 16'hff6f;
#10;
address_ina = 206;
address_inb = 207;
data_ina = 16'hfbfa;
data_inb = 16'h1cf;
#10;
address_ina = 208;
address_inb = 209;
data_ina = 16'hff3b;
data_inb = 16'hfa4e;
#10;
address_ina = 210;
address_inb = 211;
data_ina = 16'hfdf6;
data_inb = 16'hfc1f;
#10;
address_ina = 212;
address_inb = 213;
data_ina = 16'hdd;
data_inb = 16'hfe53;
#10;
address_ina = 214;
address_inb = 215;
data_ina = 16'h5f5;
data_inb = 16'h55a;
#10;
address_ina = 216;
address_inb = 217;
data_ina = 16'h18;
data_inb = 16'h150;
#10;
address_ina = 218;
address_inb = 219;
data_ina = 16'h3ac;
data_inb = 16'h284;
#10;
address_ina = 220;
address_inb = 221;
data_ina = 16'hfefb;
data_inb = 16'hfdd7;
#10;
address_ina = 222;
address_inb = 223;
data_ina = 16'hfdcd;
data_inb = 16'hfddc;
#10;
address_ina = 224;
address_inb = 225;
data_ina = 16'h59d;
data_inb = 16'hfc26;
#10;
address_ina = 226;
address_inb = 227;
data_ina = 16'hffaa;
data_inb = 16'h4ae;
#10;
address_ina = 228;
address_inb = 229;
data_ina = 16'hf9f7;
data_inb = 16'h7a;
#10;
address_ina = 230;
address_inb = 231;
data_ina = 16'hfb3d;
data_inb = 16'h4ce;
#10;
address_ina = 232;
address_inb = 233;
data_ina = 16'h52b;
data_inb = 16'h64c;
#10;
address_ina = 234;
address_inb = 235;
data_ina = 16'h40c;
data_inb = 16'h2ad;
#10;
address_ina = 236;
address_inb = 237;
data_ina = 16'h9e;
data_inb = 16'h4fe;
#10;
address_ina = 238;
address_inb = 239;
data_ina = 16'h3f3;
data_inb = 16'h271;
#10;
address_ina = 240;
address_inb = 241;
data_ina = 16'h9f;
data_inb = 16'h4d;
#10;
address_ina = 242;
address_inb = 243;
data_ina = 16'h45c;
data_inb = 16'hff42;
#10;
address_ina = 244;
address_inb = 245;
data_ina = 16'h4e4;
data_inb = 16'h2f0;
#10;
address_ina = 246;
address_inb = 247;
data_ina = 16'h5ed;
data_inb = 16'hfd3f;
#10;
address_ina = 248;
address_inb = 249;
data_ina = 16'h40b;
data_inb = 16'h372;
#10;
address_ina = 250;
address_inb = 251;
data_ina = 16'hfebe;
data_inb = 16'h174;
#10;
address_ina = 252;
address_inb = 253;
data_ina = 16'hfce5;
data_inb = 16'h33f;
#10;
address_ina = 254;
address_inb = 255;
data_ina = 16'hfc6a;
data_inb = 16'hfff9;
#10;
        wait(init_done);
        #30
        we = 0;
        // Start processing
         
		  #38000

        start = 0;



//        wait (wr_req);
//		  wait (!wr_req);
//		   rd_req = 1;
		  wait(done);
		  #20000
rd_req = 1;
        #70 
		  start = 1;
		 #80 
wait(rd_empty)
rd_req = 0;

$display("Finished the NTT test Number %d",test_num);
////Begin test number #93//////////////
rst = 1;

//#1000
start = 1;
mode = 1; //NTT 0 // INTT 1

// Reset for a few clock cycles

#1000

rst = 0;
test_num = test_num + 1;
#1000
we = 1;
address_ina = 0;
address_inb = 1;
data_ina = 16'hff62;
data_inb = 16'h125;
#10;
address_ina = 2;
address_inb = 3;
data_ina = 16'h11f;
data_inb = 16'hfc90;
#10;
address_ina = 4;
address_inb = 5;
data_ina = 16'h231;
data_inb = 16'h3d2;
#10;
address_ina = 6;
address_inb = 7;
data_ina = 16'hfdd3;
data_inb = 16'h3cd;
#10;
address_ina = 8;
address_inb = 9;
data_ina = 16'h3ef;
data_inb = 16'hcc;
#10;
address_ina = 10;
address_inb = 11;
data_ina = 16'h14;
data_inb = 16'h156;
#10;
address_ina = 12;
address_inb = 13;
data_ina = 16'h403;
data_inb = 16'h4f3;
#10;
address_ina = 14;
address_inb = 15;
data_ina = 16'h372;
data_inb = 16'h2ab;
#10;
address_ina = 16;
address_inb = 17;
data_ina = 16'h49e;
data_inb = 16'hfab5;
#10;
address_ina = 18;
address_inb = 19;
data_ina = 16'hfae0;
data_inb = 16'h593;
#10;
address_ina = 20;
address_inb = 21;
data_ina = 16'h1ac;
data_inb = 16'hfd53;
#10;
address_ina = 22;
address_inb = 23;
data_ina = 16'hfad8;
data_inb = 16'hff38;
#10;
address_ina = 24;
address_inb = 25;
data_ina = 16'hfca6;
data_inb = 16'h2a2;
#10;
address_ina = 26;
address_inb = 27;
data_ina = 16'hff76;
data_inb = 16'h4e8;
#10;
address_ina = 28;
address_inb = 29;
data_ina = 16'h680;
data_inb = 16'h309;
#10;
address_ina = 30;
address_inb = 31;
data_ina = 16'h4e5;
data_inb = 16'h5d0;
#10;
address_ina = 32;
address_inb = 33;
data_ina = 16'h113;
data_inb = 16'hff05;
#10;
address_ina = 34;
address_inb = 35;
data_ina = 16'h176;
data_inb = 16'h1f1;
#10;
address_ina = 36;
address_inb = 37;
data_ina = 16'hfe58;
data_inb = 16'h56e;
#10;
address_ina = 38;
address_inb = 39;
data_ina = 16'hfeb2;
data_inb = 16'h3f7;
#10;
address_ina = 40;
address_inb = 41;
data_ina = 16'h5cd;
data_inb = 16'h2e7;
#10;
address_ina = 42;
address_inb = 43;
data_ina = 16'hfa73;
data_inb = 16'hf9a8;
#10;
address_ina = 44;
address_inb = 45;
data_ina = 16'h60d;
data_inb = 16'hfb36;
#10;
address_ina = 46;
address_inb = 47;
data_ina = 16'h193;
data_inb = 16'h484;
#10;
address_ina = 48;
address_inb = 49;
data_ina = 16'hfd12;
data_inb = 16'hfbbe;
#10;
address_ina = 50;
address_inb = 51;
data_ina = 16'hfd69;
data_inb = 16'h42c;
#10;
address_ina = 52;
address_inb = 53;
data_ina = 16'h2b6;
data_inb = 16'hfe3b;
#10;
address_ina = 54;
address_inb = 55;
data_ina = 16'h115;
data_inb = 16'hf9d5;
#10;
address_ina = 56;
address_inb = 57;
data_ina = 16'hdd;
data_inb = 16'hf9ee;
#10;
address_ina = 58;
address_inb = 59;
data_ina = 16'h424;
data_inb = 16'hfe90;
#10;
address_ina = 60;
address_inb = 61;
data_ina = 16'h158;
data_inb = 16'hfb30;
#10;
address_ina = 62;
address_inb = 63;
data_ina = 16'h490;
data_inb = 16'hfa47;
#10;
address_ina = 64;
address_inb = 65;
data_ina = 16'h70;
data_inb = 16'h15a;
#10;
address_ina = 66;
address_inb = 67;
data_ina = 16'hfcb5;
data_inb = 16'hfd4d;
#10;
address_ina = 68;
address_inb = 69;
data_ina = 16'hfaa4;
data_inb = 16'h476;
#10;
address_ina = 70;
address_inb = 71;
data_ina = 16'hfe2d;
data_inb = 16'hfac7;
#10;
address_ina = 72;
address_inb = 73;
data_ina = 16'h119;
data_inb = 16'h527;
#10;
address_ina = 74;
address_inb = 75;
data_ina = 16'hffe3;
data_inb = 16'hfd77;
#10;
address_ina = 76;
address_inb = 77;
data_ina = 16'hfdf7;
data_inb = 16'hfd2b;
#10;
address_ina = 78;
address_inb = 79;
data_ina = 16'hfb0b;
data_inb = 16'h5fb;
#10;
address_ina = 80;
address_inb = 81;
data_ina = 16'h228;
data_inb = 16'hfbe9;
#10;
address_ina = 82;
address_inb = 83;
data_ina = 16'hfe34;
data_inb = 16'hfbc7;
#10;
address_ina = 84;
address_inb = 85;
data_ina = 16'h5b4;
data_inb = 16'hfbf3;
#10;
address_ina = 86;
address_inb = 87;
data_ina = 16'h4f8;
data_inb = 16'hfb75;
#10;
address_ina = 88;
address_inb = 89;
data_ina = 16'hfe9e;
data_inb = 16'hfe01;
#10;
address_ina = 90;
address_inb = 91;
data_ina = 16'h4bf;
data_inb = 16'h1b0;
#10;
address_ina = 92;
address_inb = 93;
data_ina = 16'h3a7;
data_inb = 16'hfd0d;
#10;
address_ina = 94;
address_inb = 95;
data_ina = 16'h623;
data_inb = 16'hfd85;
#10;
address_ina = 96;
address_inb = 97;
data_ina = 16'h3ea;
data_inb = 16'hfde7;
#10;
address_ina = 98;
address_inb = 99;
data_ina = 16'h364;
data_inb = 16'hfa9b;
#10;
address_ina = 100;
address_inb = 101;
data_ina = 16'hfc4b;
data_inb = 16'hfcaf;
#10;
address_ina = 102;
address_inb = 103;
data_ina = 16'h49a;
data_inb = 16'h66b;
#10;
address_ina = 104;
address_inb = 105;
data_ina = 16'hfcd4;
data_inb = 16'h2e2;
#10;
address_ina = 106;
address_inb = 107;
data_ina = 16'hff14;
data_inb = 16'h2d2;
#10;
address_ina = 108;
address_inb = 109;
data_ina = 16'h2a6;
data_inb = 16'h39e;
#10;
address_ina = 110;
address_inb = 111;
data_ina = 16'hfffc;
data_inb = 16'h15e;
#10;
address_ina = 112;
address_inb = 113;
data_ina = 16'h411;
data_inb = 16'hf9ec;
#10;
address_ina = 114;
address_inb = 115;
data_ina = 16'h1ac;
data_inb = 16'hffee;
#10;
address_ina = 116;
address_inb = 117;
data_ina = 16'hff19;
data_inb = 16'hfdc6;
#10;
address_ina = 118;
address_inb = 119;
data_ina = 16'hfdc8;
data_inb = 16'hdc;
#10;
address_ina = 120;
address_inb = 121;
data_ina = 16'hfc23;
data_inb = 16'hfde3;
#10;
address_ina = 122;
address_inb = 123;
data_ina = 16'h438;
data_inb = 16'hfb0a;
#10;
address_ina = 124;
address_inb = 125;
data_ina = 16'h38;
data_inb = 16'h1c3;
#10;
address_ina = 126;
address_inb = 127;
data_ina = 16'h31a;
data_inb = 16'hfe52;
#10;
address_ina = 128;
address_inb = 129;
data_ina = 16'hfbfb;
data_inb = 16'h58;
#10;
address_ina = 130;
address_inb = 131;
data_ina = 16'hfb97;
data_inb = 16'hfe3f;
#10;
address_ina = 132;
address_inb = 133;
data_ina = 16'hfa78;
data_inb = 16'hf9c6;
#10;
address_ina = 134;
address_inb = 135;
data_ina = 16'hfa46;
data_inb = 16'hfa79;
#10;
address_ina = 136;
address_inb = 137;
data_ina = 16'hfc19;
data_inb = 16'h29;
#10;
address_ina = 138;
address_inb = 139;
data_ina = 16'hfc5c;
data_inb = 16'h2d8;
#10;
address_ina = 140;
address_inb = 141;
data_ina = 16'hfda1;
data_inb = 16'h451;
#10;
address_ina = 142;
address_inb = 143;
data_ina = 16'hfde0;
data_inb = 16'hfb4a;
#10;
address_ina = 144;
address_inb = 145;
data_ina = 16'hfa81;
data_inb = 16'h5dd;
#10;
address_ina = 146;
address_inb = 147;
data_ina = 16'h5a4;
data_inb = 16'hfdaf;
#10;
address_ina = 148;
address_inb = 149;
data_ina = 16'hf9f8;
data_inb = 16'h3a3;
#10;
address_ina = 150;
address_inb = 151;
data_ina = 16'hff11;
data_inb = 16'hfa65;
#10;
address_ina = 152;
address_inb = 153;
data_ina = 16'hff16;
data_inb = 16'h4f0;
#10;
address_ina = 154;
address_inb = 155;
data_ina = 16'hfdce;
data_inb = 16'h668;
#10;
address_ina = 156;
address_inb = 157;
data_ina = 16'h311;
data_inb = 16'h168;
#10;
address_ina = 158;
address_inb = 159;
data_ina = 16'hfe8a;
data_inb = 16'hfa91;
#10;
address_ina = 160;
address_inb = 161;
data_ina = 16'hfa99;
data_inb = 16'h578;
#10;
address_ina = 162;
address_inb = 163;
data_ina = 16'h234;
data_inb = 16'hfb99;
#10;
address_ina = 164;
address_inb = 165;
data_ina = 16'h3c4;
data_inb = 16'h1df;
#10;
address_ina = 166;
address_inb = 167;
data_ina = 16'hff80;
data_inb = 16'h31c;
#10;
address_ina = 168;
address_inb = 169;
data_ina = 16'hfba2;
data_inb = 16'hfb44;
#10;
address_ina = 170;
address_inb = 171;
data_ina = 16'h3ca;
data_inb = 16'hfb1a;
#10;
address_ina = 172;
address_inb = 173;
data_ina = 16'h570;
data_inb = 16'h3d4;
#10;
address_ina = 174;
address_inb = 175;
data_ina = 16'hfd33;
data_inb = 16'h3e;
#10;
address_ina = 176;
address_inb = 177;
data_ina = 16'hfed2;
data_inb = 16'hfddc;
#10;
address_ina = 178;
address_inb = 179;
data_ina = 16'hfecb;
data_inb = 16'hfe93;
#10;
address_ina = 180;
address_inb = 181;
data_ina = 16'hfb29;
data_inb = 16'hfbbc;
#10;
address_ina = 182;
address_inb = 183;
data_ina = 16'hf9e4;
data_inb = 16'hfc1a;
#10;
address_ina = 184;
address_inb = 185;
data_ina = 16'hfb9d;
data_inb = 16'h40e;
#10;
address_ina = 186;
address_inb = 187;
data_ina = 16'h2c2;
data_inb = 16'hfe36;
#10;
address_ina = 188;
address_inb = 189;
data_ina = 16'h2;
data_inb = 16'hfe84;
#10;
address_ina = 190;
address_inb = 191;
data_ina = 16'hfb64;
data_inb = 16'h567;
#10;
address_ina = 192;
address_inb = 193;
data_ina = 16'h1d5;
data_inb = 16'h3bc;
#10;
address_ina = 194;
address_inb = 195;
data_ina = 16'h652;
data_inb = 16'hfa0d;
#10;
address_ina = 196;
address_inb = 197;
data_ina = 16'h40b;
data_inb = 16'hff23;
#10;
address_ina = 198;
address_inb = 199;
data_ina = 16'h14d;
data_inb = 16'h205;
#10;
address_ina = 200;
address_inb = 201;
data_ina = 16'hfab7;
data_inb = 16'hf98c;
#10;
address_ina = 202;
address_inb = 203;
data_ina = 16'hfe4d;
data_inb = 16'hfe5e;
#10;
address_ina = 204;
address_inb = 205;
data_ina = 16'h4a0;
data_inb = 16'hfe60;
#10;
address_ina = 206;
address_inb = 207;
data_ina = 16'h427;
data_inb = 16'hfa1a;
#10;
address_ina = 208;
address_inb = 209;
data_ina = 16'hfb39;
data_inb = 16'h173;
#10;
address_ina = 210;
address_inb = 211;
data_ina = 16'hcb;
data_inb = 16'h5cb;
#10;
address_ina = 212;
address_inb = 213;
data_ina = 16'h34b;
data_inb = 16'h2b7;
#10;
address_ina = 214;
address_inb = 215;
data_ina = 16'h31e;
data_inb = 16'hfe87;
#10;
address_ina = 216;
address_inb = 217;
data_ina = 16'h48b;
data_inb = 16'hfb2f;
#10;
address_ina = 218;
address_inb = 219;
data_ina = 16'hfe8e;
data_inb = 16'hff5e;
#10;
address_ina = 220;
address_inb = 221;
data_ina = 16'h2f7;
data_inb = 16'h327;
#10;
address_ina = 222;
address_inb = 223;
data_ina = 16'h561;
data_inb = 16'hfa76;
#10;
address_ina = 224;
address_inb = 225;
data_ina = 16'hfaa1;
data_inb = 16'h20d;
#10;
address_ina = 226;
address_inb = 227;
data_ina = 16'h4cf;
data_inb = 16'h175;
#10;
address_ina = 228;
address_inb = 229;
data_ina = 16'h3a;
data_inb = 16'hf9d7;
#10;
address_ina = 230;
address_inb = 231;
data_ina = 16'hfef1;
data_inb = 16'hfd17;
#10;
address_ina = 232;
address_inb = 233;
data_ina = 16'h1e8;
data_inb = 16'h23e;
#10;
address_ina = 234;
address_inb = 235;
data_ina = 16'hfdd4;
data_inb = 16'h527;
#10;
address_ina = 236;
address_inb = 237;
data_ina = 16'h615;
data_inb = 16'hf9b0;
#10;
address_ina = 238;
address_inb = 239;
data_ina = 16'h580;
data_inb = 16'h44b;
#10;
address_ina = 240;
address_inb = 241;
data_ina = 16'hfac6;
data_inb = 16'h96;
#10;
address_ina = 242;
address_inb = 243;
data_ina = 16'hff8a;
data_inb = 16'hfcb6;
#10;
address_ina = 244;
address_inb = 245;
data_ina = 16'hfe68;
data_inb = 16'h21e;
#10;
address_ina = 246;
address_inb = 247;
data_ina = 16'hfdc0;
data_inb = 16'h2c1;
#10;
address_ina = 248;
address_inb = 249;
data_ina = 16'hfd0d;
data_inb = 16'hfaba;
#10;
address_ina = 250;
address_inb = 251;
data_ina = 16'h1a6;
data_inb = 16'hfcca;
#10;
address_ina = 252;
address_inb = 253;
data_ina = 16'hfd2e;
data_inb = 16'h57;
#10;
address_ina = 254;
address_inb = 255;
data_ina = 16'hfb7c;
data_inb = 16'hfea5;
#10;
        wait(init_done);
        #30
        we = 0;
        // Start processing
         
		  #38000

        start = 0;



//        wait (wr_req);
//		  wait (!wr_req);
//		   rd_req = 1;
		  wait(done);
		  #20000
rd_req = 1;
        #70 
		  start = 1;
		 #80 
wait(rd_empty)
rd_req = 0;

$display("Finished the NTT test Number %d",test_num);
////Begin test number #94//////////////
rst = 1;

//#1000
start = 1;
mode = 0; //NTT 0 // INTT 1

// Reset for a few clock cycles

#1000

rst = 0;
test_num = test_num + 1;
#1000
we = 1;
address_ina = 0;
address_inb = 1;
data_ina = 16'hce7;
data_inb = 16'h80d;
#10;
address_ina = 2;
address_inb = 3;
data_ina = 16'h4b0;
data_inb = 16'ha2c;
#10;
address_ina = 4;
address_inb = 5;
data_ina = 16'h2a;
data_inb = 16'h145;
#10;
address_ina = 6;
address_inb = 7;
data_ina = 16'h837;
data_inb = 16'h74d;
#10;
address_ina = 8;
address_inb = 9;
data_ina = 16'h55f;
data_inb = 16'h504;
#10;
address_ina = 10;
address_inb = 11;
data_ina = 16'h3ac;
data_inb = 16'h8ea;
#10;
address_ina = 12;
address_inb = 13;
data_ina = 16'h7a8;
data_inb = 16'h96;
#10;
address_ina = 14;
address_inb = 15;
data_ina = 16'h236;
data_inb = 16'h8c0;
#10;
address_ina = 16;
address_inb = 17;
data_ina = 16'h4ed;
data_inb = 16'ha70;
#10;
address_ina = 18;
address_inb = 19;
data_ina = 16'h9fb;
data_inb = 16'hb40;
#10;
address_ina = 20;
address_inb = 21;
data_ina = 16'h13b;
data_inb = 16'h28a;
#10;
address_ina = 22;
address_inb = 23;
data_ina = 16'h979;
data_inb = 16'hcb3;
#10;
address_ina = 24;
address_inb = 25;
data_ina = 16'haa4;
data_inb = 16'h85e;
#10;
address_ina = 26;
address_inb = 27;
data_ina = 16'hc48;
data_inb = 16'ha81;
#10;
address_ina = 28;
address_inb = 29;
data_ina = 16'h774;
data_inb = 16'hb09;
#10;
address_ina = 30;
address_inb = 31;
data_ina = 16'h1bd;
data_inb = 16'h9eb;
#10;
address_ina = 32;
address_inb = 33;
data_ina = 16'h525;
data_inb = 16'h11e;
#10;
address_ina = 34;
address_inb = 35;
data_ina = 16'h89f;
data_inb = 16'h13b;
#10;
address_ina = 36;
address_inb = 37;
data_ina = 16'h785;
data_inb = 16'h78;
#10;
address_ina = 38;
address_inb = 39;
data_ina = 16'h2d5;
data_inb = 16'h8bd;
#10;
address_ina = 40;
address_inb = 41;
data_ina = 16'h80a;
data_inb = 16'h5c4;
#10;
address_ina = 42;
address_inb = 43;
data_ina = 16'h62c;
data_inb = 16'h323;
#10;
address_ina = 44;
address_inb = 45;
data_ina = 16'h6dc;
data_inb = 16'h899;
#10;
address_ina = 46;
address_inb = 47;
data_ina = 16'hbd3;
data_inb = 16'h5e4;
#10;
address_ina = 48;
address_inb = 49;
data_ina = 16'h53b;
data_inb = 16'hb2a;
#10;
address_ina = 50;
address_inb = 51;
data_ina = 16'ha60;
data_inb = 16'h538;
#10;
address_ina = 52;
address_inb = 53;
data_ina = 16'hfe;
data_inb = 16'h10b;
#10;
address_ina = 54;
address_inb = 55;
data_ina = 16'h6a8;
data_inb = 16'h63f;
#10;
address_ina = 56;
address_inb = 57;
data_ina = 16'h86f;
data_inb = 16'hc3;
#10;
address_ina = 58;
address_inb = 59;
data_ina = 16'hb7e;
data_inb = 16'hbcc;
#10;
address_ina = 60;
address_inb = 61;
data_ina = 16'h421;
data_inb = 16'h284;
#10;
address_ina = 62;
address_inb = 63;
data_ina = 16'h96c;
data_inb = 16'h3;
#10;
address_ina = 64;
address_inb = 65;
data_ina = 16'h336;
data_inb = 16'h989;
#10;
address_ina = 66;
address_inb = 67;
data_ina = 16'haf6;
data_inb = 16'h1c7;
#10;
address_ina = 68;
address_inb = 69;
data_ina = 16'hac5;
data_inb = 16'h53f;
#10;
address_ina = 70;
address_inb = 71;
data_ina = 16'h367;
data_inb = 16'haa8;
#10;
address_ina = 72;
address_inb = 73;
data_ina = 16'h569;
data_inb = 16'h2e8;
#10;
address_ina = 74;
address_inb = 75;
data_ina = 16'h6e2;
data_inb = 16'h166;
#10;
address_ina = 76;
address_inb = 77;
data_ina = 16'h344;
data_inb = 16'h5e;
#10;
address_ina = 78;
address_inb = 79;
data_ina = 16'h918;
data_inb = 16'h844;
#10;
address_ina = 80;
address_inb = 81;
data_ina = 16'h218;
data_inb = 16'h27;
#10;
address_ina = 82;
address_inb = 83;
data_ina = 16'h807;
data_inb = 16'h444;
#10;
address_ina = 84;
address_inb = 85;
data_ina = 16'h13f;
data_inb = 16'hc9c;
#10;
address_ina = 86;
address_inb = 87;
data_ina = 16'ha77;
data_inb = 16'h703;
#10;
address_ina = 88;
address_inb = 89;
data_ina = 16'h92;
data_inb = 16'hb2d;
#10;
address_ina = 90;
address_inb = 91;
data_ina = 16'h907;
data_inb = 16'hce4;
#10;
address_ina = 92;
address_inb = 93;
data_ina = 16'h5ce;
data_inb = 16'h19a;
#10;
address_ina = 94;
address_inb = 95;
data_ina = 16'h64c;
data_inb = 16'hab5;
#10;
address_ina = 96;
address_inb = 97;
data_ina = 16'h663;
data_inb = 16'hae5;
#10;
address_ina = 98;
address_inb = 99;
data_ina = 16'h973;
data_inb = 16'h44;
#10;
address_ina = 100;
address_inb = 101;
data_ina = 16'h576;
data_inb = 16'h458;
#10;
address_ina = 102;
address_inb = 103;
data_ina = 16'h5ee;
data_inb = 16'h5a0;
#10;
address_ina = 104;
address_inb = 105;
data_ina = 16'h569;
data_inb = 16'h824;
#10;
address_ina = 106;
address_inb = 107;
data_ina = 16'ha05;
data_inb = 16'haf9;
#10;
address_ina = 108;
address_inb = 109;
data_ina = 16'hb6;
data_inb = 16'h9aa;
#10;
address_ina = 110;
address_inb = 111;
data_ina = 16'hbfa;
data_inb = 16'h485;
#10;
address_ina = 112;
address_inb = 113;
data_ina = 16'h205;
data_inb = 16'h2c5;
#10;
address_ina = 114;
address_inb = 115;
data_ina = 16'h3f3;
data_inb = 16'hab1;
#10;
address_ina = 116;
address_inb = 117;
data_ina = 16'ha3;
data_inb = 16'hbfa;
#10;
address_ina = 118;
address_inb = 119;
data_ina = 16'h525;
data_inb = 16'h441;
#10;
address_ina = 120;
address_inb = 121;
data_ina = 16'hc21;
data_inb = 16'h5ba;
#10;
address_ina = 122;
address_inb = 123;
data_ina = 16'h441;
data_inb = 16'h8b6;
#10;
address_ina = 124;
address_inb = 125;
data_ina = 16'h28d;
data_inb = 16'h3f3;
#10;
address_ina = 126;
address_inb = 127;
data_ina = 16'h9cb;
data_inb = 16'h40d;
#10;
address_ina = 128;
address_inb = 129;
data_ina = 16'h2f9;
data_inb = 16'h663;
#10;
address_ina = 130;
address_inb = 131;
data_ina = 16'h4b9;
data_inb = 16'haf2;
#10;
address_ina = 132;
address_inb = 133;
data_ina = 16'hcc0;
data_inb = 16'h45b;
#10;
address_ina = 134;
address_inb = 135;
data_ina = 16'h62f;
data_inb = 16'h344;
#10;
address_ina = 136;
address_inb = 137;
data_ina = 16'h3a5;
data_inb = 16'h7c6;
#10;
address_ina = 138;
address_inb = 139;
data_ina = 16'h3d6;
data_inb = 16'h50e;
#10;
address_ina = 140;
address_inb = 141;
data_ina = 16'h280;
data_inb = 16'h521;
#10;
address_ina = 142;
address_inb = 143;
data_ina = 16'ha6d;
data_inb = 16'ha50;
#10;
address_ina = 144;
address_inb = 145;
data_ina = 16'h36e;
data_inb = 16'hb0c;
#10;
address_ina = 146;
address_inb = 147;
data_ina = 16'h2b4;
data_inb = 16'he0;
#10;
address_ina = 148;
address_inb = 149;
data_ina = 16'hced;
data_inb = 16'h378;
#10;
address_ina = 150;
address_inb = 151;
data_ina = 16'h5b0;
data_inb = 16'h3b5;
#10;
address_ina = 152;
address_inb = 153;
data_ina = 16'h196;
data_inb = 16'h458;
#10;
address_ina = 154;
address_inb = 155;
data_ina = 16'h5b;
data_inb = 16'h7bc;
#10;
address_ina = 156;
address_inb = 157;
data_ina = 16'h34d;
data_inb = 16'hca;
#10;
address_ina = 158;
address_inb = 159;
data_ina = 16'h107;
data_inb = 16'h4bd;
#10;
address_ina = 160;
address_inb = 161;
data_ina = 16'h107;
data_inb = 16'h2f2;
#10;
address_ina = 162;
address_inb = 163;
data_ina = 16'h4cd;
data_inb = 16'hc96;
#10;
address_ina = 164;
address_inb = 165;
data_ina = 16'ha5a;
data_inb = 16'h202;
#10;
address_ina = 166;
address_inb = 167;
data_ina = 16'h15c;
data_inb = 16'h61c;
#10;
address_ina = 168;
address_inb = 169;
data_ina = 16'h266;
data_inb = 16'h74a;
#10;
address_ina = 170;
address_inb = 171;
data_ina = 16'h4e0;
data_inb = 16'h4f7;
#10;
address_ina = 172;
address_inb = 173;
data_ina = 16'h945;
data_inb = 16'h663;
#10;
address_ina = 174;
address_inb = 175;
data_ina = 16'h639;
data_inb = 16'h650;
#10;
address_ina = 176;
address_inb = 177;
data_ina = 16'h465;
data_inb = 16'h166;
#10;
address_ina = 178;
address_inb = 179;
data_ina = 16'h93b;
data_inb = 16'h9f2;
#10;
address_ina = 180;
address_inb = 181;
data_ina = 16'hc17;
data_inb = 16'h865;
#10;
address_ina = 182;
address_inb = 183;
data_ina = 16'he0;
data_inb = 16'h1a;
#10;
address_ina = 184;
address_inb = 185;
data_ina = 16'hcdd;
data_inb = 16'h3ac;
#10;
address_ina = 186;
address_inb = 187;
data_ina = 16'h6b5;
data_inb = 16'h434;
#10;
address_ina = 188;
address_inb = 189;
data_ina = 16'hcb9;
data_inb = 16'h589;
#10;
address_ina = 190;
address_inb = 191;
data_ina = 16'ha33;
data_inb = 16'h79f;
#10;
address_ina = 192;
address_inb = 193;
data_ina = 16'h414;
data_inb = 16'h20f;
#10;
address_ina = 194;
address_inb = 195;
data_ina = 16'h6ec;
data_inb = 16'h38e;
#10;
address_ina = 196;
address_inb = 197;
data_ina = 16'h4a6;
data_inb = 16'h8e7;
#10;
address_ina = 198;
address_inb = 199;
data_ina = 16'haab;
data_inb = 16'h11e;
#10;
address_ina = 200;
address_inb = 201;
data_ina = 16'h403;
data_inb = 16'h848;
#10;
address_ina = 202;
address_inb = 203;
data_ina = 16'h666;
data_inb = 16'h42e;
#10;
address_ina = 204;
address_inb = 205;
data_ina = 16'h62;
data_inb = 16'hbbf;
#10;
address_ina = 206;
address_inb = 207;
data_ina = 16'h414;
data_inb = 16'h107;
#10;
address_ina = 208;
address_inb = 209;
data_ina = 16'h4c0;
data_inb = 16'h43b;
#10;
address_ina = 210;
address_inb = 211;
data_ina = 16'h18d;
data_inb = 16'hb4d;
#10;
address_ina = 212;
address_inb = 213;
data_ina = 16'ha84;
data_inb = 16'h670;
#10;
address_ina = 214;
address_inb = 215;
data_ina = 16'h6b1;
data_inb = 16'h455;
#10;
address_ina = 216;
address_inb = 217;
data_ina = 16'h55;
data_inb = 16'h6dc;
#10;
address_ina = 218;
address_inb = 219;
data_ina = 16'ha77;
data_inb = 16'hac5;
#10;
address_ina = 220;
address_inb = 221;
data_ina = 16'h10e;
data_inb = 16'h11e;
#10;
address_ina = 222;
address_inb = 223;
data_ina = 16'h3a5;
data_inb = 16'h3b;
#10;
address_ina = 224;
address_inb = 225;
data_ina = 16'h6c8;
data_inb = 16'hc72;
#10;
address_ina = 226;
address_inb = 227;
data_ina = 16'haf9;
data_inb = 16'hbb9;
#10;
address_ina = 228;
address_inb = 229;
data_ina = 16'h9d1;
data_inb = 16'h302;
#10;
address_ina = 230;
address_inb = 231;
data_ina = 16'ha9b;
data_inb = 16'hc4e;
#10;
address_ina = 232;
address_inb = 233;
data_ina = 16'h1d7;
data_inb = 16'h65d;
#10;
address_ina = 234;
address_inb = 235;
data_ina = 16'hc44;
data_inb = 16'hc3;
#10;
address_ina = 236;
address_inb = 237;
data_ina = 16'h552;
data_inb = 16'hcf4;
#10;
address_ina = 238;
address_inb = 239;
data_ina = 16'h3d3;
data_inb = 16'h8f;
#10;
address_ina = 240;
address_inb = 241;
data_ina = 16'h9e8;
data_inb = 16'h1c1;
#10;
address_ina = 242;
address_inb = 243;
data_ina = 16'h798;
data_inb = 16'h485;
#10;
address_ina = 244;
address_inb = 245;
data_ina = 16'h6bb;
data_inb = 16'hced;
#10;
address_ina = 246;
address_inb = 247;
data_ina = 16'hc2e;
data_inb = 16'h6dc;
#10;
address_ina = 248;
address_inb = 249;
data_ina = 16'h5a3;
data_inb = 16'h663;
#10;
address_ina = 250;
address_inb = 251;
data_ina = 16'h875;
data_inb = 16'h821;
#10;
address_ina = 252;
address_inb = 253;
data_ina = 16'ha60;
data_inb = 16'h8ed;
#10;
address_ina = 254;
address_inb = 255;
data_ina = 16'h60b;
data_inb = 16'h3dc;
#10;
        wait(init_done);
        #30
        we = 0;
        // Start processing
         
		  #38000

        start = 0;



//        wait (wr_req);
//		  wait (!wr_req);
//		   rd_req = 1;
		  wait(done);
		  #20000
rd_req = 1;
        #70 
		  start = 1;
		 #80 
wait(rd_empty)
rd_req = 0;

$display("Finished the NTT test Number %d",test_num);
////Begin test number #95//////////////
rst = 1;

//#1000
start = 1;
mode = 0; //NTT 0 // INTT 1

// Reset for a few clock cycles

#1000

rst = 0;
test_num = test_num + 1;
#1000
we = 1;
address_ina = 0;
address_inb = 1;
data_ina = 16'h817;
data_inb = 16'hc1a;
#10;
address_ina = 2;
address_inb = 3;
data_ina = 16'h378;
data_inb = 16'h1bd;
#10;
address_ina = 4;
address_inb = 5;
data_ina = 16'hb74;
data_inb = 16'h525;
#10;
address_ina = 6;
address_inb = 7;
data_ina = 16'h4b6;
data_inb = 16'h28d;
#10;
address_ina = 8;
address_inb = 9;
data_ina = 16'h7d3;
data_inb = 16'h2b8;
#10;
address_ina = 10;
address_inb = 11;
data_ina = 16'hfe;
data_inb = 16'h7bc;
#10;
address_ina = 12;
address_inb = 13;
data_ina = 16'h5fb;
data_inb = 16'haa8;
#10;
address_ina = 14;
address_inb = 15;
data_ina = 16'h99a;
data_inb = 16'ha0f;
#10;
address_ina = 16;
address_inb = 17;
data_ina = 16'h2a;
data_inb = 16'h1d;
#10;
address_ina = 18;
address_inb = 19;
data_ina = 16'h3e;
data_inb = 16'h1ad;
#10;
address_ina = 20;
address_inb = 21;
data_ina = 16'h246;
data_inb = 16'h580;
#10;
address_ina = 22;
address_inb = 23;
data_ina = 16'h3b5;
data_inb = 16'h67a;
#10;
address_ina = 24;
address_inb = 25;
data_ina = 16'hbb5;
data_inb = 16'h499;
#10;
address_ina = 26;
address_inb = 27;
data_ina = 16'h104;
data_inb = 16'h6e5;
#10;
address_ina = 28;
address_inb = 29;
data_ina = 16'h1b0;
data_inb = 16'h761;
#10;
address_ina = 30;
address_inb = 31;
data_ina = 16'h3b2;
data_inb = 16'h193;
#10;
address_ina = 32;
address_inb = 33;
data_ina = 16'h482;
data_inb = 16'h79f;
#10;
address_ina = 34;
address_inb = 35;
data_ina = 16'h1a7;
data_inb = 16'h444;
#10;
address_ina = 36;
address_inb = 37;
data_ina = 16'h1f1;
data_inb = 16'h10b;
#10;
address_ina = 38;
address_inb = 39;
data_ina = 16'ha4d;
data_inb = 16'h367;
#10;
address_ina = 40;
address_inb = 41;
data_ina = 16'h525;
data_inb = 16'h5ba;
#10;
address_ina = 42;
address_inb = 43;
data_ina = 16'hc41;
data_inb = 16'h347;
#10;
address_ina = 44;
address_inb = 45;
data_ina = 16'h858;
data_inb = 16'h542;
#10;
address_ina = 46;
address_inb = 47;
data_ina = 16'h277;
data_inb = 16'hab5;
#10;
address_ina = 48;
address_inb = 49;
data_ina = 16'h589;
data_inb = 16'h68e;
#10;
address_ina = 50;
address_inb = 51;
data_ina = 16'h1c4;
data_inb = 16'h65d;
#10;
address_ina = 52;
address_inb = 53;
data_ina = 16'h6f2;
data_inb = 16'h733;
#10;
address_ina = 54;
address_inb = 55;
data_ina = 16'ha26;
data_inb = 16'hb74;
#10;
address_ina = 56;
address_inb = 57;
data_ina = 16'h8c3;
data_inb = 16'h911;
#10;
address_ina = 58;
address_inb = 59;
data_ina = 16'h67d;
data_inb = 16'hbd;
#10;
address_ina = 60;
address_inb = 61;
data_ina = 16'h8e0;
data_inb = 16'h85b;
#10;
address_ina = 62;
address_inb = 63;
data_ina = 16'h9a3;
data_inb = 16'h2ce;
#10;
address_ina = 64;
address_inb = 65;
data_ina = 16'h23f;
data_inb = 16'ha5d;
#10;
address_ina = 66;
address_inb = 67;
data_ina = 16'h653;
data_inb = 16'h1d4;
#10;
address_ina = 68;
address_inb = 69;
data_ina = 16'hb40;
data_inb = 16'h5eb;
#10;
address_ina = 70;
address_inb = 71;
data_ina = 16'h2d2;
data_inb = 16'hbd;
#10;
address_ina = 72;
address_inb = 73;
data_ina = 16'hbfa;
data_inb = 16'hc37;
#10;
address_ina = 74;
address_inb = 75;
data_ina = 16'h673;
data_inb = 16'h9cb;
#10;
address_ina = 76;
address_inb = 77;
data_ina = 16'h2ce;
data_inb = 16'haf6;
#10;
address_ina = 78;
address_inb = 79;
data_ina = 16'h68a;
data_inb = 16'h3c6;
#10;
address_ina = 80;
address_inb = 81;
data_ina = 16'h7af;
data_inb = 16'hb6b;
#10;
address_ina = 82;
address_inb = 83;
data_ina = 16'h5f1;
data_inb = 16'h8ed;
#10;
address_ina = 84;
address_inb = 85;
data_ina = 16'h90b;
data_inb = 16'h7e3;
#10;
address_ina = 86;
address_inb = 87;
data_ina = 16'h111;
data_inb = 16'hb8b;
#10;
address_ina = 88;
address_inb = 89;
data_ina = 16'h489;
data_inb = 16'h7fa;
#10;
address_ina = 90;
address_inb = 91;
data_ina = 16'h757;
data_inb = 16'h1c1;
#10;
address_ina = 92;
address_inb = 93;
data_ina = 16'h3b;
data_inb = 16'h7dc;
#10;
address_ina = 94;
address_inb = 95;
data_ina = 16'h284;
data_inb = 16'hb06;
#10;
address_ina = 96;
address_inb = 97;
data_ina = 16'hb81;
data_inb = 16'h911;
#10;
address_ina = 98;
address_inb = 99;
data_ina = 16'h3bf;
data_inb = 16'h455;
#10;
address_ina = 100;
address_inb = 101;
data_ina = 16'hcc3;
data_inb = 16'hbe9;
#10;
address_ina = 102;
address_inb = 103;
data_ina = 16'ha26;
data_inb = 16'h138;
#10;
address_ina = 104;
address_inb = 105;
data_ina = 16'h3d9;
data_inb = 16'h618;
#10;
address_ina = 106;
address_inb = 107;
data_ina = 16'h5f5;
data_inb = 16'h1b4;
#10;
address_ina = 108;
address_inb = 109;
data_ina = 16'h20f;
data_inb = 16'h94f;
#10;
address_ina = 110;
address_inb = 111;
data_ina = 16'h99;
data_inb = 16'h834;
#10;
address_ina = 112;
address_inb = 113;
data_ina = 16'h159;
data_inb = 16'ha5a;
#10;
address_ina = 114;
address_inb = 115;
data_ina = 16'hb7e;
data_inb = 16'h7ac;
#10;
address_ina = 116;
address_inb = 117;
data_ina = 16'h63c;
data_inb = 16'h8a3;
#10;
address_ina = 118;
address_inb = 119;
data_ina = 16'h179;
data_inb = 16'h3af;
#10;
address_ina = 120;
address_inb = 121;
data_ina = 16'h8fe;
data_inb = 16'h111;
#10;
address_ina = 122;
address_inb = 123;
data_ina = 16'h9ff;
data_inb = 16'h740;
#10;
address_ina = 124;
address_inb = 125;
data_ina = 16'h212;
data_inb = 16'h284;
#10;
address_ina = 126;
address_inb = 127;
data_ina = 16'h22c;
data_inb = 16'hcd3;
#10;
address_ina = 128;
address_inb = 129;
data_ina = 16'h189;
data_inb = 16'h492;
#10;
address_ina = 130;
address_inb = 131;
data_ina = 16'h9f8;
data_inb = 16'h253;
#10;
address_ina = 132;
address_inb = 133;
data_ina = 16'h5ca;
data_inb = 16'h918;
#10;
address_ina = 134;
address_inb = 135;
data_ina = 16'h159;
data_inb = 16'h485;
#10;
address_ina = 136;
address_inb = 137;
data_ina = 16'h618;
data_inb = 16'h55c;
#10;
address_ina = 138;
address_inb = 139;
data_ina = 16'h2ff;
data_inb = 16'ha08;
#10;
address_ina = 140;
address_inb = 141;
data_ina = 16'hc44;
data_inb = 16'h5fb;
#10;
address_ina = 142;
address_inb = 143;
data_ina = 16'hc92;
data_inb = 16'h966;
#10;
address_ina = 144;
address_inb = 145;
data_ina = 16'hca6;
data_inb = 16'h521;
#10;
address_ina = 146;
address_inb = 147;
data_ina = 16'h5d7;
data_inb = 16'hba8;
#10;
address_ina = 148;
address_inb = 149;
data_ina = 16'h844;
data_inb = 16'h72d;
#10;
address_ina = 150;
address_inb = 151;
data_ina = 16'ha2c;
data_inb = 16'h684;
#10;
address_ina = 152;
address_inb = 153;
data_ina = 16'h99;
data_inb = 16'h41a;
#10;
address_ina = 154;
address_inb = 155;
data_ina = 16'h1ad;
data_inb = 16'h8e0;
#10;
address_ina = 156;
address_inb = 157;
data_ina = 16'h26d;
data_inb = 16'h17;
#10;
address_ina = 158;
address_inb = 159;
data_ina = 16'h733;
data_inb = 16'hb4a;
#10;
address_ina = 160;
address_inb = 161;
data_ina = 16'h417;
data_inb = 16'h96f;
#10;
address_ina = 162;
address_inb = 163;
data_ina = 16'h81a;
data_inb = 16'h3af;
#10;
address_ina = 164;
address_inb = 165;
data_ina = 16'h27a;
data_inb = 16'h54f;
#10;
address_ina = 166;
address_inb = 167;
data_ina = 16'h7;
data_inb = 16'h407;
#10;
address_ina = 168;
address_inb = 169;
data_ina = 16'h2c5;
data_inb = 16'hbd6;
#10;
address_ina = 170;
address_inb = 171;
data_ina = 16'h7c;
data_inb = 16'h649;
#10;
address_ina = 172;
address_inb = 173;
data_ina = 16'hd7;
data_inb = 16'ha05;
#10;
address_ina = 174;
address_inb = 175;
data_ina = 16'h7af;
data_inb = 16'hc48;
#10;
address_ina = 176;
address_inb = 177;
data_ina = 16'h583;
data_inb = 16'h74a;
#10;
address_ina = 178;
address_inb = 179;
data_ina = 16'hc41;
data_inb = 16'h885;
#10;
address_ina = 180;
address_inb = 181;
data_ina = 16'h754;
data_inb = 16'hc14;
#10;
address_ina = 182;
address_inb = 183;
data_ina = 16'h61f;
data_inb = 16'h3fd;
#10;
address_ina = 184;
address_inb = 185;
data_ina = 16'h9b0;
data_inb = 16'h973;
#10;
address_ina = 186;
address_inb = 187;
data_ina = 16'ha5d;
data_inb = 16'h29a;
#10;
address_ina = 188;
address_inb = 189;
data_ina = 16'h8d0;
data_inb = 16'h761;
#10;
address_ina = 190;
address_inb = 191;
data_ina = 16'h417;
data_inb = 16'h7b9;
#10;
address_ina = 192;
address_inb = 193;
data_ina = 16'h9bd;
data_inb = 16'h266;
#10;
address_ina = 194;
address_inb = 195;
data_ina = 16'hc6f;
data_inb = 16'h896;
#10;
address_ina = 196;
address_inb = 197;
data_ina = 16'h82a;
data_inb = 16'h173;
#10;
address_ina = 198;
address_inb = 199;
data_ina = 16'hc3b;
data_inb = 16'ha4d;
#10;
address_ina = 200;
address_inb = 201;
data_ina = 16'h3d6;
data_inb = 16'h9e8;
#10;
address_ina = 202;
address_inb = 203;
data_ina = 16'h593;
data_inb = 16'h8a3;
#10;
address_ina = 204;
address_inb = 205;
data_ina = 16'ha84;
data_inb = 16'h225;
#10;
address_ina = 206;
address_inb = 207;
data_ina = 16'h605;
data_inb = 16'h6bb;
#10;
address_ina = 208;
address_inb = 209;
data_ina = 16'hc55;
data_inb = 16'h6f;
#10;
address_ina = 210;
address_inb = 211;
data_ina = 16'h8ac;
data_inb = 16'h448;
#10;
address_ina = 212;
address_inb = 213;
data_ina = 16'h79f;
data_inb = 16'h6a1;
#10;
address_ina = 214;
address_inb = 215;
data_ina = 16'h1b4;
data_inb = 16'hba5;
#10;
address_ina = 216;
address_inb = 217;
data_ina = 16'h7b5;
data_inb = 16'hcc0;
#10;
address_ina = 218;
address_inb = 219;
data_ina = 16'h4b0;
data_inb = 16'hc62;
#10;
address_ina = 220;
address_inb = 221;
data_ina = 16'h72d;
data_inb = 16'h831;
#10;
address_ina = 222;
address_inb = 223;
data_ina = 16'h7a8;
data_inb = 16'haa8;
#10;
address_ina = 224;
address_inb = 225;
data_ina = 16'h173;
data_inb = 16'haef;
#10;
address_ina = 226;
address_inb = 227;
data_ina = 16'h326;
data_inb = 16'h4b;
#10;
address_ina = 228;
address_inb = 229;
data_ina = 16'hb03;
data_inb = 16'h778;
#10;
address_ina = 230;
address_inb = 231;
data_ina = 16'hf1;
data_inb = 16'h7a5;
#10;
address_ina = 232;
address_inb = 233;
data_ina = 16'h1b7;
data_inb = 16'h169;
#10;
address_ina = 234;
address_inb = 235;
data_ina = 16'h7cc;
data_inb = 16'h78;
#10;
address_ina = 236;
address_inb = 237;
data_ina = 16'h9cb;
data_inb = 16'h2df;
#10;
address_ina = 238;
address_inb = 239;
data_ina = 16'h1b4;
data_inb = 16'hc3;
#10;
address_ina = 240;
address_inb = 241;
data_ina = 16'h848;
data_inb = 16'hbf6;
#10;
address_ina = 242;
address_inb = 243;
data_ina = 16'ha8e;
data_inb = 16'h492;
#10;
address_ina = 244;
address_inb = 245;
data_ina = 16'h431;
data_inb = 16'h6ef;
#10;
address_ina = 246;
address_inb = 247;
data_ina = 16'hfe;
data_inb = 16'h361;
#10;
address_ina = 248;
address_inb = 249;
data_ina = 16'h928;
data_inb = 16'h932;
#10;
address_ina = 250;
address_inb = 251;
data_ina = 16'h499;
data_inb = 16'hc9f;
#10;
address_ina = 252;
address_inb = 253;
data_ina = 16'ha7d;
data_inb = 16'h2b1;
#10;
address_ina = 254;
address_inb = 255;
data_ina = 16'hb2a;
data_inb = 16'h5de;
#10;
        wait(init_done);
        #30
        we = 0;
        // Start processing
         
		  #38000

        start = 0;



//        wait (wr_req);
//		  wait (!wr_req);
//		   rd_req = 1;
		  wait(done);
		  #20000
rd_req = 1;
        #70 
		  start = 1;
		 #80 
wait(rd_empty)
rd_req = 0;

$display("Finished the NTT test Number %d",test_num);
////Begin test number #96//////////////
rst = 1;

//#1000
start = 1;
mode = 1; //NTT 0 // INTT 1

// Reset for a few clock cycles

#1000

rst = 0;
test_num = test_num + 1;
#1000
we = 1;
address_ina = 0;
address_inb = 1;
data_ina = 16'hcc;
data_inb = 16'hfa4b;
#10;
address_ina = 2;
address_inb = 3;
data_ina = 16'hfa01;
data_inb = 16'h4c6;
#10;
address_ina = 4;
address_inb = 5;
data_ina = 16'hfb6f;
data_inb = 16'hfc64;
#10;
address_ina = 6;
address_inb = 7;
data_ina = 16'h495;
data_inb = 16'hfff1;
#10;
address_ina = 8;
address_inb = 9;
data_ina = 16'hff9c;
data_inb = 16'hfc73;
#10;
address_ina = 10;
address_inb = 11;
data_ina = 16'h203;
data_inb = 16'hfc34;
#10;
address_ina = 12;
address_inb = 13;
data_ina = 16'hfcd6;
data_inb = 16'h567;
#10;
address_ina = 14;
address_inb = 15;
data_ina = 16'h301;
data_inb = 16'h19b;
#10;
address_ina = 16;
address_inb = 17;
data_ina = 16'h327;
data_inb = 16'h471;
#10;
address_ina = 18;
address_inb = 19;
data_ina = 16'hfd8c;
data_inb = 16'h1e8;
#10;
address_ina = 20;
address_inb = 21;
data_ina = 16'h450;
data_inb = 16'hff96;
#10;
address_ina = 22;
address_inb = 23;
data_ina = 16'h2c1;
data_inb = 16'hfb83;
#10;
address_ina = 24;
address_inb = 25;
data_ina = 16'h292;
data_inb = 16'hfe64;
#10;
address_ina = 26;
address_inb = 27;
data_ina = 16'hffb2;
data_inb = 16'h499;
#10;
address_ina = 28;
address_inb = 29;
data_ina = 16'hc3;
data_inb = 16'hfa08;
#10;
address_ina = 30;
address_inb = 31;
data_ina = 16'hfa39;
data_inb = 16'hfdda;
#10;
address_ina = 32;
address_inb = 33;
data_ina = 16'h4e;
data_inb = 16'hfaee;
#10;
address_ina = 34;
address_inb = 35;
data_ina = 16'hfdec;
data_inb = 16'h3ed;
#10;
address_ina = 36;
address_inb = 37;
data_ina = 16'hfd97;
data_inb = 16'hfe14;
#10;
address_ina = 38;
address_inb = 39;
data_ina = 16'h11c;
data_inb = 16'hfcc6;
#10;
address_ina = 40;
address_inb = 41;
data_ina = 16'hed;
data_inb = 16'hfa83;
#10;
address_ina = 42;
address_inb = 43;
data_ina = 16'hff56;
data_inb = 16'h47a;
#10;
address_ina = 44;
address_inb = 45;
data_ina = 16'h1e1;
data_inb = 16'h606;
#10;
address_ina = 46;
address_inb = 47;
data_ina = 16'hfcf4;
data_inb = 16'hfbc2;
#10;
address_ina = 48;
address_inb = 49;
data_ina = 16'hfb15;
data_inb = 16'hfbe9;
#10;
address_ina = 50;
address_inb = 51;
data_ina = 16'h202;
data_inb = 16'h346;
#10;
address_ina = 52;
address_inb = 53;
data_ina = 16'h218;
data_inb = 16'hfcc8;
#10;
address_ina = 54;
address_inb = 55;
data_ina = 16'h329;
data_inb = 16'hfe97;
#10;
address_ina = 56;
address_inb = 57;
data_ina = 16'hfa88;
data_inb = 16'h145;
#10;
address_ina = 58;
address_inb = 59;
data_ina = 16'h45f;
data_inb = 16'h4e0;
#10;
address_ina = 60;
address_inb = 61;
data_ina = 16'h3cf;
data_inb = 16'hff23;
#10;
address_ina = 62;
address_inb = 63;
data_ina = 16'h517;
data_inb = 16'h454;
#10;
address_ina = 64;
address_inb = 65;
data_ina = 16'h29b;
data_inb = 16'h65b;
#10;
address_ina = 66;
address_inb = 67;
data_ina = 16'hfaac;
data_inb = 16'hfe96;
#10;
address_ina = 68;
address_inb = 69;
data_ina = 16'hff77;
data_inb = 16'hfff2;
#10;
address_ina = 70;
address_inb = 71;
data_ina = 16'hff15;
data_inb = 16'h5fc;
#10;
address_ina = 72;
address_inb = 73;
data_ina = 16'hfeba;
data_inb = 16'h59a;
#10;
address_ina = 74;
address_inb = 75;
data_ina = 16'h3c4;
data_inb = 16'hfccb;
#10;
address_ina = 76;
address_inb = 77;
data_ina = 16'h15c;
data_inb = 16'hfa5e;
#10;
address_ina = 78;
address_inb = 79;
data_ina = 16'hd0;
data_inb = 16'h430;
#10;
address_ina = 80;
address_inb = 81;
data_ina = 16'h3a3;
data_inb = 16'h76;
#10;
address_ina = 82;
address_inb = 83;
data_ina = 16'hffa7;
data_inb = 16'hff33;
#10;
address_ina = 84;
address_inb = 85;
data_ina = 16'hfc3a;
data_inb = 16'h54e;
#10;
address_ina = 86;
address_inb = 87;
data_ina = 16'h49f;
data_inb = 16'hfca4;
#10;
address_ina = 88;
address_inb = 89;
data_ina = 16'h2ac;
data_inb = 16'h63c;
#10;
address_ina = 90;
address_inb = 91;
data_ina = 16'h46c;
data_inb = 16'hfc32;
#10;
address_ina = 92;
address_inb = 93;
data_ina = 16'h1ba;
data_inb = 16'h504;
#10;
address_ina = 94;
address_inb = 95;
data_ina = 16'hfcf8;
data_inb = 16'h76;
#10;
address_ina = 96;
address_inb = 97;
data_ina = 16'hfeba;
data_inb = 16'h5ea;
#10;
address_ina = 98;
address_inb = 99;
data_ina = 16'h3f1;
data_inb = 16'h2cd;
#10;
address_ina = 100;
address_inb = 101;
data_ina = 16'hfc31;
data_inb = 16'hfe4b;
#10;
address_ina = 102;
address_inb = 103;
data_ina = 16'h5e9;
data_inb = 16'h7d;
#10;
address_ina = 104;
address_inb = 105;
data_ina = 16'hfd3f;
data_inb = 16'hfbd8;
#10;
address_ina = 106;
address_inb = 107;
data_ina = 16'h2be;
data_inb = 16'h561;
#10;
address_ina = 108;
address_inb = 109;
data_ina = 16'h57f;
data_inb = 16'h5a4;
#10;
address_ina = 110;
address_inb = 111;
data_ina = 16'h61a;
data_inb = 16'h41e;
#10;
address_ina = 112;
address_inb = 113;
data_ina = 16'h4ef;
data_inb = 16'hfa33;
#10;
address_ina = 114;
address_inb = 115;
data_ina = 16'he7;
data_inb = 16'hfa92;
#10;
address_ina = 116;
address_inb = 117;
data_ina = 16'h5a6;
data_inb = 16'h416;
#10;
address_ina = 118;
address_inb = 119;
data_ina = 16'h4d7;
data_inb = 16'hfb83;
#10;
address_ina = 120;
address_inb = 121;
data_ina = 16'hff70;
data_inb = 16'hfffb;
#10;
address_ina = 122;
address_inb = 123;
data_ina = 16'hfba7;
data_inb = 16'hfa94;
#10;
address_ina = 124;
address_inb = 125;
data_ina = 16'h5a6;
data_inb = 16'h25f;
#10;
address_ina = 126;
address_inb = 127;
data_ina = 16'h30a;
data_inb = 16'h27a;
#10;
address_ina = 128;
address_inb = 129;
data_ina = 16'hfdea;
data_inb = 16'hfbed;
#10;
address_ina = 130;
address_inb = 131;
data_ina = 16'hfaab;
data_inb = 16'h3e0;
#10;
address_ina = 132;
address_inb = 133;
data_ina = 16'hfc11;
data_inb = 16'hfc91;
#10;
address_ina = 134;
address_inb = 135;
data_ina = 16'hfcc6;
data_inb = 16'h329;
#10;
address_ina = 136;
address_inb = 137;
data_ina = 16'hfa20;
data_inb = 16'h605;
#10;
address_ina = 138;
address_inb = 139;
data_ina = 16'h25e;
data_inb = 16'h114;
#10;
address_ina = 140;
address_inb = 141;
data_ina = 16'h304;
data_inb = 16'h396;
#10;
address_ina = 142;
address_inb = 143;
data_ina = 16'hfd1f;
data_inb = 16'hac;
#10;
address_ina = 144;
address_inb = 145;
data_ina = 16'hfde0;
data_inb = 16'hfd33;
#10;
address_ina = 146;
address_inb = 147;
data_ina = 16'h454;
data_inb = 16'hfe2a;
#10;
address_ina = 148;
address_inb = 149;
data_ina = 16'h5f;
data_inb = 16'h5c9;
#10;
address_ina = 150;
address_inb = 151;
data_ina = 16'hfdd9;
data_inb = 16'hfd15;
#10;
address_ina = 152;
address_inb = 153;
data_ina = 16'hffc3;
data_inb = 16'hfbf9;
#10;
address_ina = 154;
address_inb = 155;
data_ina = 16'hfca5;
data_inb = 16'hff6d;
#10;
address_ina = 156;
address_inb = 157;
data_ina = 16'h40d;
data_inb = 16'h176;
#10;
address_ina = 158;
address_inb = 159;
data_ina = 16'h523;
data_inb = 16'h522;
#10;
address_ina = 160;
address_inb = 161;
data_ina = 16'hfe54;
data_inb = 16'h27;
#10;
address_ina = 162;
address_inb = 163;
data_ina = 16'hfb7c;
data_inb = 16'hfecc;
#10;
address_ina = 164;
address_inb = 165;
data_ina = 16'h1c0;
data_inb = 16'h500;
#10;
address_ina = 166;
address_inb = 167;
data_ina = 16'hfa96;
data_inb = 16'h2f0;
#10;
address_ina = 168;
address_inb = 169;
data_ina = 16'hfcde;
data_inb = 16'hfa9d;
#10;
address_ina = 170;
address_inb = 171;
data_ina = 16'h277;
data_inb = 16'hfbb2;
#10;
address_ina = 172;
address_inb = 173;
data_ina = 16'h341;
data_inb = 16'h680;
#10;
address_ina = 174;
address_inb = 175;
data_ina = 16'h66;
data_inb = 16'h663;
#10;
address_ina = 176;
address_inb = 177;
data_ina = 16'h65c;
data_inb = 16'h401;
#10;
address_ina = 178;
address_inb = 179;
data_ina = 16'h4e9;
data_inb = 16'hfab8;
#10;
address_ina = 180;
address_inb = 181;
data_ina = 16'hfe64;
data_inb = 16'hfa0f;
#10;
address_ina = 182;
address_inb = 183;
data_ina = 16'h1f1;
data_inb = 16'hfdea;
#10;
address_ina = 184;
address_inb = 185;
data_ina = 16'hfbb9;
data_inb = 16'h321;
#10;
address_ina = 186;
address_inb = 187;
data_ina = 16'h2ef;
data_inb = 16'hfa93;
#10;
address_ina = 188;
address_inb = 189;
data_ina = 16'hfbe4;
data_inb = 16'hfeab;
#10;
address_ina = 190;
address_inb = 191;
data_ina = 16'h295;
data_inb = 16'h22f;
#10;
address_ina = 192;
address_inb = 193;
data_ina = 16'hfdf9;
data_inb = 16'hfa6a;
#10;
address_ina = 194;
address_inb = 195;
data_ina = 16'h3f8;
data_inb = 16'h679;
#10;
address_ina = 196;
address_inb = 197;
data_ina = 16'hfa67;
data_inb = 16'h17;
#10;
address_ina = 198;
address_inb = 199;
data_ina = 16'h13;
data_inb = 16'h3de;
#10;
address_ina = 200;
address_inb = 201;
data_ina = 16'hfcb7;
data_inb = 16'hfd20;
#10;
address_ina = 202;
address_inb = 203;
data_ina = 16'hfa60;
data_inb = 16'h436;
#10;
address_ina = 204;
address_inb = 205;
data_ina = 16'h3c9;
data_inb = 16'hfe06;
#10;
address_ina = 206;
address_inb = 207;
data_ina = 16'h379;
data_inb = 16'h58a;
#10;
address_ina = 208;
address_inb = 209;
data_ina = 16'hff53;
data_inb = 16'h58b;
#10;
address_ina = 210;
address_inb = 211;
data_ina = 16'hff2b;
data_inb = 16'hfdf2;
#10;
address_ina = 212;
address_inb = 213;
data_ina = 16'hfd00;
data_inb = 16'hfa7e;
#10;
address_ina = 214;
address_inb = 215;
data_ina = 16'h3fd;
data_inb = 16'hff1a;
#10;
address_ina = 216;
address_inb = 217;
data_ina = 16'hfbcd;
data_inb = 16'hfaa5;
#10;
address_ina = 218;
address_inb = 219;
data_ina = 16'hfdf9;
data_inb = 16'h139;
#10;
address_ina = 220;
address_inb = 221;
data_ina = 16'h41e;
data_inb = 16'hf9cf;
#10;
address_ina = 222;
address_inb = 223;
data_ina = 16'h5d;
data_inb = 16'hfac1;
#10;
address_ina = 224;
address_inb = 225;
data_ina = 16'hfdba;
data_inb = 16'h244;
#10;
address_ina = 226;
address_inb = 227;
data_ina = 16'h13e;
data_inb = 16'h521;
#10;
address_ina = 228;
address_inb = 229;
data_ina = 16'h491;
data_inb = 16'hffa4;
#10;
address_ina = 230;
address_inb = 231;
data_ina = 16'h539;
data_inb = 16'hf9ed;
#10;
address_ina = 232;
address_inb = 233;
data_ina = 16'h522;
data_inb = 16'h1a6;
#10;
address_ina = 234;
address_inb = 235;
data_ina = 16'h3c0;
data_inb = 16'hfd53;
#10;
address_ina = 236;
address_inb = 237;
data_ina = 16'h66d;
data_inb = 16'hfa41;
#10;
address_ina = 238;
address_inb = 239;
data_ina = 16'hf9a5;
data_inb = 16'hfb7f;
#10;
address_ina = 240;
address_inb = 241;
data_ina = 16'he6;
data_inb = 16'hfb30;
#10;
address_ina = 242;
address_inb = 243;
data_ina = 16'hfaea;
data_inb = 16'h33a;
#10;
address_ina = 244;
address_inb = 245;
data_ina = 16'h3b5;
data_inb = 16'hfdb9;
#10;
address_ina = 246;
address_inb = 247;
data_ina = 16'h241;
data_inb = 16'h4f5;
#10;
address_ina = 248;
address_inb = 249;
data_ina = 16'hfbb5;
data_inb = 16'hfdea;
#10;
address_ina = 250;
address_inb = 251;
data_ina = 16'h578;
data_inb = 16'h464;
#10;
address_ina = 252;
address_inb = 253;
data_ina = 16'hfdee;
data_inb = 16'hff38;
#10;
address_ina = 254;
address_inb = 255;
data_ina = 16'hfa91;
data_inb = 16'h634;
#10;
        wait(init_done);
        #30
        we = 0;
        // Start processing
         
		  #38000

        start = 0;



//        wait (wr_req);
//		  wait (!wr_req);
//		   rd_req = 1;
		  wait(done);
		  #20000
rd_req = 1;
        #70 
		  start = 1;
		 #80 
wait(rd_empty)
rd_req = 0;

$display("Finished the NTT test Number %d",test_num);
////Begin test number #97//////////////
rst = 1;

//#1000
start = 1;
mode = 0; //NTT 0 // INTT 1

// Reset for a few clock cycles

#1000

rst = 0;
test_num = test_num + 1;
#1000
we = 1;
address_ina = 0;
address_inb = 1;
data_ina = 16'hffff;
data_inb = 16'h3;
#10;
address_ina = 2;
address_inb = 3;
data_ina = 16'h0;
data_inb = 16'hfffe;
#10;
address_ina = 4;
address_inb = 5;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 6;
address_inb = 7;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 8;
address_inb = 9;
data_ina = 16'hffff;
data_inb = 16'h2;
#10;
address_ina = 10;
address_inb = 11;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 12;
address_inb = 13;
data_ina = 16'h2;
data_inb = 16'h0;
#10;
address_ina = 14;
address_inb = 15;
data_ina = 16'h2;
data_inb = 16'hfffe;
#10;
address_ina = 16;
address_inb = 17;
data_ina = 16'hfffe;
data_inb = 16'h2;
#10;
address_ina = 18;
address_inb = 19;
data_ina = 16'hfffd;
data_inb = 16'hffff;
#10;
address_ina = 20;
address_inb = 21;
data_ina = 16'h3;
data_inb = 16'h0;
#10;
address_ina = 22;
address_inb = 23;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 24;
address_inb = 25;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 26;
address_inb = 27;
data_ina = 16'h0;
data_inb = 16'h3;
#10;
address_ina = 28;
address_inb = 29;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 30;
address_inb = 31;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 32;
address_inb = 33;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 34;
address_inb = 35;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 36;
address_inb = 37;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 38;
address_inb = 39;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 40;
address_inb = 41;
data_ina = 16'hfffe;
data_inb = 16'hffff;
#10;
address_ina = 42;
address_inb = 43;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 44;
address_inb = 45;
data_ina = 16'hffff;
data_inb = 16'h2;
#10;
address_ina = 46;
address_inb = 47;
data_ina = 16'hfffd;
data_inb = 16'h0;
#10;
address_ina = 48;
address_inb = 49;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 50;
address_inb = 51;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 52;
address_inb = 53;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 54;
address_inb = 55;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 56;
address_inb = 57;
data_ina = 16'hfffe;
data_inb = 16'hffff;
#10;
address_ina = 58;
address_inb = 59;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 60;
address_inb = 61;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 62;
address_inb = 63;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 64;
address_inb = 65;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 66;
address_inb = 67;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 68;
address_inb = 69;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 70;
address_inb = 71;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 72;
address_inb = 73;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 74;
address_inb = 75;
data_ina = 16'h2;
data_inb = 16'h1;
#10;
address_ina = 76;
address_inb = 77;
data_ina = 16'h0;
data_inb = 16'h2;
#10;
address_ina = 78;
address_inb = 79;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 80;
address_inb = 81;
data_ina = 16'h1;
data_inb = 16'hfffe;
#10;
address_ina = 82;
address_inb = 83;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 84;
address_inb = 85;
data_ina = 16'hffff;
data_inb = 16'hfffe;
#10;
address_ina = 86;
address_inb = 87;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 88;
address_inb = 89;
data_ina = 16'h0;
data_inb = 16'hfffe;
#10;
address_ina = 90;
address_inb = 91;
data_ina = 16'h2;
data_inb = 16'h0;
#10;
address_ina = 92;
address_inb = 93;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 94;
address_inb = 95;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 96;
address_inb = 97;
data_ina = 16'hfffe;
data_inb = 16'h2;
#10;
address_ina = 98;
address_inb = 99;
data_ina = 16'hfffe;
data_inb = 16'h1;
#10;
address_ina = 100;
address_inb = 101;
data_ina = 16'h0;
data_inb = 16'h2;
#10;
address_ina = 102;
address_inb = 103;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 104;
address_inb = 105;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 106;
address_inb = 107;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 108;
address_inb = 109;
data_ina = 16'h1;
data_inb = 16'hfffe;
#10;
address_ina = 110;
address_inb = 111;
data_ina = 16'hfffe;
data_inb = 16'hffff;
#10;
address_ina = 112;
address_inb = 113;
data_ina = 16'hfffe;
data_inb = 16'h1;
#10;
address_ina = 114;
address_inb = 115;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 116;
address_inb = 117;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 118;
address_inb = 119;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 120;
address_inb = 121;
data_ina = 16'h2;
data_inb = 16'hfffd;
#10;
address_ina = 122;
address_inb = 123;
data_ina = 16'h2;
data_inb = 16'hfffe;
#10;
address_ina = 124;
address_inb = 125;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 126;
address_inb = 127;
data_ina = 16'h1;
data_inb = 16'hfffd;
#10;
address_ina = 128;
address_inb = 129;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 130;
address_inb = 131;
data_ina = 16'h2;
data_inb = 16'hfffe;
#10;
address_ina = 132;
address_inb = 133;
data_ina = 16'h2;
data_inb = 16'h0;
#10;
address_ina = 134;
address_inb = 135;
data_ina = 16'h2;
data_inb = 16'hfffe;
#10;
address_ina = 136;
address_inb = 137;
data_ina = 16'h0;
data_inb = 16'h2;
#10;
address_ina = 138;
address_inb = 139;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 140;
address_inb = 141;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 142;
address_inb = 143;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 144;
address_inb = 145;
data_ina = 16'h2;
data_inb = 16'hfffe;
#10;
address_ina = 146;
address_inb = 147;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 148;
address_inb = 149;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 150;
address_inb = 151;
data_ina = 16'h2;
data_inb = 16'h1;
#10;
address_ina = 152;
address_inb = 153;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 154;
address_inb = 155;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 156;
address_inb = 157;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 158;
address_inb = 159;
data_ina = 16'h1;
data_inb = 16'hfffe;
#10;
address_ina = 160;
address_inb = 161;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 162;
address_inb = 163;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 164;
address_inb = 165;
data_ina = 16'hffff;
data_inb = 16'h2;
#10;
address_ina = 166;
address_inb = 167;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 168;
address_inb = 169;
data_ina = 16'h3;
data_inb = 16'h0;
#10;
address_ina = 170;
address_inb = 171;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 172;
address_inb = 173;
data_ina = 16'hffff;
data_inb = 16'hfffe;
#10;
address_ina = 174;
address_inb = 175;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 176;
address_inb = 177;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 178;
address_inb = 179;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 180;
address_inb = 181;
data_ina = 16'h2;
data_inb = 16'h1;
#10;
address_ina = 182;
address_inb = 183;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 184;
address_inb = 185;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 186;
address_inb = 187;
data_ina = 16'h0;
data_inb = 16'h3;
#10;
address_ina = 188;
address_inb = 189;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 190;
address_inb = 191;
data_ina = 16'h0;
data_inb = 16'hfffe;
#10;
address_ina = 192;
address_inb = 193;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 194;
address_inb = 195;
data_ina = 16'h0;
data_inb = 16'hfffe;
#10;
address_ina = 196;
address_inb = 197;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 198;
address_inb = 199;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 200;
address_inb = 201;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 202;
address_inb = 203;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 204;
address_inb = 205;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 206;
address_inb = 207;
data_ina = 16'h1;
data_inb = 16'hfffe;
#10;
address_ina = 208;
address_inb = 209;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 210;
address_inb = 211;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 212;
address_inb = 213;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 214;
address_inb = 215;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 216;
address_inb = 217;
data_ina = 16'hffff;
data_inb = 16'hfffd;
#10;
address_ina = 218;
address_inb = 219;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 220;
address_inb = 221;
data_ina = 16'h0;
data_inb = 16'h2;
#10;
address_ina = 222;
address_inb = 223;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 224;
address_inb = 225;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 226;
address_inb = 227;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 228;
address_inb = 229;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 230;
address_inb = 231;
data_ina = 16'h2;
data_inb = 16'h1;
#10;
address_ina = 232;
address_inb = 233;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 234;
address_inb = 235;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 236;
address_inb = 237;
data_ina = 16'h2;
data_inb = 16'h2;
#10;
address_ina = 238;
address_inb = 239;
data_ina = 16'h3;
data_inb = 16'h0;
#10;
address_ina = 240;
address_inb = 241;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 242;
address_inb = 243;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 244;
address_inb = 245;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 246;
address_inb = 247;
data_ina = 16'h2;
data_inb = 16'h1;
#10;
address_ina = 248;
address_inb = 249;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 250;
address_inb = 251;
data_ina = 16'h0;
data_inb = 16'hfffe;
#10;
address_ina = 252;
address_inb = 253;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 254;
address_inb = 255;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
        wait(init_done);
        #30
        we = 0;
        // Start processing
         
		  #38000

        start = 0;



//        wait (wr_req);
//		  wait (!wr_req);
//		   rd_req = 1;
		  wait(done);
		  #20000
rd_req = 1;
        #70 
		  start = 1;
		 #80 
wait(rd_empty)
rd_req = 0;

$display("Finished the NTT test Number %d",test_num);
////Begin test number #98//////////////
rst = 1;

//#1000
start = 1;
mode = 0; //NTT 0 // INTT 1

// Reset for a few clock cycles

#1000

rst = 0;
test_num = test_num + 1;
#1000
we = 1;
address_ina = 0;
address_inb = 1;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 2;
address_inb = 3;
data_ina = 16'h2;
data_inb = 16'h0;
#10;
address_ina = 4;
address_inb = 5;
data_ina = 16'hffff;
data_inb = 16'h2;
#10;
address_ina = 6;
address_inb = 7;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 8;
address_inb = 9;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 10;
address_inb = 11;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 12;
address_inb = 13;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 14;
address_inb = 15;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 16;
address_inb = 17;
data_ina = 16'h0;
data_inb = 16'h2;
#10;
address_ina = 18;
address_inb = 19;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 20;
address_inb = 21;
data_ina = 16'hfffe;
data_inb = 16'h0;
#10;
address_ina = 22;
address_inb = 23;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 24;
address_inb = 25;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 26;
address_inb = 27;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 28;
address_inb = 29;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 30;
address_inb = 31;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 32;
address_inb = 33;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 34;
address_inb = 35;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 36;
address_inb = 37;
data_ina = 16'h2;
data_inb = 16'hfffe;
#10;
address_ina = 38;
address_inb = 39;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 40;
address_inb = 41;
data_ina = 16'h1;
data_inb = 16'hfffe;
#10;
address_ina = 42;
address_inb = 43;
data_ina = 16'hffff;
data_inb = 16'h2;
#10;
address_ina = 44;
address_inb = 45;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 46;
address_inb = 47;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 48;
address_inb = 49;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 50;
address_inb = 51;
data_ina = 16'hfffd;
data_inb = 16'h1;
#10;
address_ina = 52;
address_inb = 53;
data_ina = 16'hfffe;
data_inb = 16'hffff;
#10;
address_ina = 54;
address_inb = 55;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 56;
address_inb = 57;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 58;
address_inb = 59;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 60;
address_inb = 61;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 62;
address_inb = 63;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 64;
address_inb = 65;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 66;
address_inb = 67;
data_ina = 16'hfffe;
data_inb = 16'hfffe;
#10;
address_ina = 68;
address_inb = 69;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 70;
address_inb = 71;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 72;
address_inb = 73;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 74;
address_inb = 75;
data_ina = 16'hfffe;
data_inb = 16'hffff;
#10;
address_ina = 76;
address_inb = 77;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 78;
address_inb = 79;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 80;
address_inb = 81;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 82;
address_inb = 83;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 84;
address_inb = 85;
data_ina = 16'hfffe;
data_inb = 16'h1;
#10;
address_ina = 86;
address_inb = 87;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 88;
address_inb = 89;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 90;
address_inb = 91;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 92;
address_inb = 93;
data_ina = 16'h0;
data_inb = 16'h2;
#10;
address_ina = 94;
address_inb = 95;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 96;
address_inb = 97;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 98;
address_inb = 99;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 100;
address_inb = 101;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 102;
address_inb = 103;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 104;
address_inb = 105;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 106;
address_inb = 107;
data_ina = 16'h2;
data_inb = 16'h0;
#10;
address_ina = 108;
address_inb = 109;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 110;
address_inb = 111;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 112;
address_inb = 113;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 114;
address_inb = 115;
data_ina = 16'h2;
data_inb = 16'h0;
#10;
address_ina = 116;
address_inb = 117;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 118;
address_inb = 119;
data_ina = 16'h3;
data_inb = 16'h3;
#10;
address_ina = 120;
address_inb = 121;
data_ina = 16'hffff;
data_inb = 16'h2;
#10;
address_ina = 122;
address_inb = 123;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 124;
address_inb = 125;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 126;
address_inb = 127;
data_ina = 16'h0;
data_inb = 16'h2;
#10;
address_ina = 128;
address_inb = 129;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 130;
address_inb = 131;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 132;
address_inb = 133;
data_ina = 16'h2;
data_inb = 16'h0;
#10;
address_ina = 134;
address_inb = 135;
data_ina = 16'h2;
data_inb = 16'hffff;
#10;
address_ina = 136;
address_inb = 137;
data_ina = 16'h0;
data_inb = 16'h3;
#10;
address_ina = 138;
address_inb = 139;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 140;
address_inb = 141;
data_ina = 16'h2;
data_inb = 16'h1;
#10;
address_ina = 142;
address_inb = 143;
data_ina = 16'h0;
data_inb = 16'hfffe;
#10;
address_ina = 144;
address_inb = 145;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 146;
address_inb = 147;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 148;
address_inb = 149;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 150;
address_inb = 151;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 152;
address_inb = 153;
data_ina = 16'h0;
data_inb = 16'hffff;
#10;
address_ina = 154;
address_inb = 155;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 156;
address_inb = 157;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 158;
address_inb = 159;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 160;
address_inb = 161;
data_ina = 16'h2;
data_inb = 16'h0;
#10;
address_ina = 162;
address_inb = 163;
data_ina = 16'h2;
data_inb = 16'hffff;
#10;
address_ina = 164;
address_inb = 165;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 166;
address_inb = 167;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 168;
address_inb = 169;
data_ina = 16'hffff;
data_inb = 16'hfffe;
#10;
address_ina = 170;
address_inb = 171;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 172;
address_inb = 173;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 174;
address_inb = 175;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 176;
address_inb = 177;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 178;
address_inb = 179;
data_ina = 16'hfffe;
data_inb = 16'h2;
#10;
address_ina = 180;
address_inb = 181;
data_ina = 16'h2;
data_inb = 16'h0;
#10;
address_ina = 182;
address_inb = 183;
data_ina = 16'h0;
data_inb = 16'hfffe;
#10;
address_ina = 184;
address_inb = 185;
data_ina = 16'h3;
data_inb = 16'h1;
#10;
address_ina = 186;
address_inb = 187;
data_ina = 16'h2;
data_inb = 16'h0;
#10;
address_ina = 188;
address_inb = 189;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 190;
address_inb = 191;
data_ina = 16'h2;
data_inb = 16'h2;
#10;
address_ina = 192;
address_inb = 193;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 194;
address_inb = 195;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 196;
address_inb = 197;
data_ina = 16'h0;
data_inb = 16'hfffe;
#10;
address_ina = 198;
address_inb = 199;
data_ina = 16'h1;
data_inb = 16'h2;
#10;
address_ina = 200;
address_inb = 201;
data_ina = 16'h0;
data_inb = 16'hfffd;
#10;
address_ina = 202;
address_inb = 203;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 204;
address_inb = 205;
data_ina = 16'h0;
data_inb = 16'h1;
#10;
address_ina = 206;
address_inb = 207;
data_ina = 16'h2;
data_inb = 16'hfffe;
#10;
address_ina = 208;
address_inb = 209;
data_ina = 16'hfffe;
data_inb = 16'h0;
#10;
address_ina = 210;
address_inb = 211;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 212;
address_inb = 213;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 214;
address_inb = 215;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 216;
address_inb = 217;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 218;
address_inb = 219;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 220;
address_inb = 221;
data_ina = 16'h2;
data_inb = 16'h0;
#10;
address_ina = 222;
address_inb = 223;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 224;
address_inb = 225;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 226;
address_inb = 227;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 228;
address_inb = 229;
data_ina = 16'hffff;
data_inb = 16'h3;
#10;
address_ina = 230;
address_inb = 231;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 232;
address_inb = 233;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
address_ina = 234;
address_inb = 235;
data_ina = 16'h1;
data_inb = 16'hffff;
#10;
address_ina = 236;
address_inb = 237;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 238;
address_inb = 239;
data_ina = 16'hfffe;
data_inb = 16'h1;
#10;
address_ina = 240;
address_inb = 241;
data_ina = 16'hffff;
data_inb = 16'hfffe;
#10;
address_ina = 242;
address_inb = 243;
data_ina = 16'h0;
data_inb = 16'h2;
#10;
address_ina = 244;
address_inb = 245;
data_ina = 16'hffff;
data_inb = 16'hffff;
#10;
address_ina = 246;
address_inb = 247;
data_ina = 16'hffff;
data_inb = 16'h1;
#10;
address_ina = 248;
address_inb = 249;
data_ina = 16'h1;
data_inb = 16'h0;
#10;
address_ina = 250;
address_inb = 251;
data_ina = 16'hffff;
data_inb = 16'h0;
#10;
address_ina = 252;
address_inb = 253;
data_ina = 16'h0;
data_inb = 16'h0;
#10;
address_ina = 254;
address_inb = 255;
data_ina = 16'h1;
data_inb = 16'h1;
#10;
        wait(init_done);
        #30
        we = 0;
        // Start processing
         
		  #38000

        start = 0;



//        wait (wr_req);
//		  wait (!wr_req);
//		   rd_req = 1;
		  wait(done);
		  #20000
rd_req = 1;
        #70 
		  start = 1;
		 #80 
wait(rd_empty)
rd_req = 0;

$display("Finished the NTT test Number %d",test_num);
////Begin test number #99//////////////
rst = 1;

//#1000
start = 1;
mode = 1; //NTT 0 // INTT 1

// Reset for a few clock cycles

#1000

rst = 0;
test_num = test_num + 1;
#1000
we = 1;
address_ina = 0;
address_inb = 1;
data_ina = 16'hfc93;
data_inb = 16'h491;
#10;
address_ina = 2;
address_inb = 3;
data_ina = 16'hfb32;
data_inb = 16'h591;
#10;
address_ina = 4;
address_inb = 5;
data_ina = 16'hfc5b;
data_inb = 16'h31c;
#10;
address_ina = 6;
address_inb = 7;
data_ina = 16'h341;
data_inb = 16'hfd3a;
#10;
address_ina = 8;
address_inb = 9;
data_ina = 16'hfbe2;
data_inb = 16'hff46;
#10;
address_ina = 10;
address_inb = 11;
data_ina = 16'hff93;
data_inb = 16'h672;
#10;
address_ina = 12;
address_inb = 13;
data_ina = 16'h34b;
data_inb = 16'hfba5;
#10;
address_ina = 14;
address_inb = 15;
data_ina = 16'h4da;
data_inb = 16'hff05;
#10;
address_ina = 16;
address_inb = 17;
data_ina = 16'h498;
data_inb = 16'hfe53;
#10;
address_ina = 18;
address_inb = 19;
data_ina = 16'hfc2b;
data_inb = 16'h62e;
#10;
address_ina = 20;
address_inb = 21;
data_ina = 16'h37c;
data_inb = 16'h603;
#10;
address_ina = 22;
address_inb = 23;
data_ina = 16'hfad8;
data_inb = 16'h654;
#10;
address_ina = 24;
address_inb = 25;
data_ina = 16'hfef1;
data_inb = 16'h593;
#10;
address_ina = 26;
address_inb = 27;
data_ina = 16'hff7e;
data_inb = 16'h4c3;
#10;
address_ina = 28;
address_inb = 29;
data_ina = 16'h324;
data_inb = 16'hfead;
#10;
address_ina = 30;
address_inb = 31;
data_ina = 16'h2b7;
data_inb = 16'hfd85;
#10;
address_ina = 32;
address_inb = 33;
data_ina = 16'h2d2;
data_inb = 16'h53d;
#10;
address_ina = 34;
address_inb = 35;
data_ina = 16'hfd45;
data_inb = 16'h3a7;
#10;
address_ina = 36;
address_inb = 37;
data_ina = 16'h35c;
data_inb = 16'hfadb;
#10;
address_ina = 38;
address_inb = 39;
data_ina = 16'hfd11;
data_inb = 16'hfe59;
#10;
address_ina = 40;
address_inb = 41;
data_ina = 16'h429;
data_inb = 16'hf986;
#10;
address_ina = 42;
address_inb = 43;
data_ina = 16'hfbb0;
data_inb = 16'hffa0;
#10;
address_ina = 44;
address_inb = 45;
data_ina = 16'hf9ab;
data_inb = 16'h306;
#10;
address_ina = 46;
address_inb = 47;
data_ina = 16'h671;
data_inb = 16'hfc0b;
#10;
address_ina = 48;
address_inb = 49;
data_ina = 16'h199;
data_inb = 16'hfcfc;
#10;
address_ina = 50;
address_inb = 51;
data_ina = 16'h605;
data_inb = 16'hff41;
#10;
address_ina = 52;
address_inb = 53;
data_ina = 16'h442;
data_inb = 16'hfa23;
#10;
address_ina = 54;
address_inb = 55;
data_ina = 16'hfb5b;
data_inb = 16'h674;
#10;
address_ina = 56;
address_inb = 57;
data_ina = 16'h2de;
data_inb = 16'h51c;
#10;
address_ina = 58;
address_inb = 59;
data_ina = 16'h7c;
data_inb = 16'h651;
#10;
address_ina = 60;
address_inb = 61;
data_ina = 16'hfd1c;
data_inb = 16'hff5a;
#10;
address_ina = 62;
address_inb = 63;
data_ina = 16'h21a;
data_inb = 16'h40c;
#10;
address_ina = 64;
address_inb = 65;
data_ina = 16'hfd43;
data_inb = 16'hfa59;
#10;
address_ina = 66;
address_inb = 67;
data_ina = 16'hfb22;
data_inb = 16'h5fa;
#10;
address_ina = 68;
address_inb = 69;
data_ina = 16'hfcab;
data_inb = 16'hfb09;
#10;
address_ina = 70;
address_inb = 71;
data_ina = 16'hffc3;
data_inb = 16'hfad1;
#10;
address_ina = 72;
address_inb = 73;
data_ina = 16'hfb74;
data_inb = 16'h63;
#10;
address_ina = 74;
address_inb = 75;
data_ina = 16'h3de;
data_inb = 16'h82;
#10;
address_ina = 76;
address_inb = 77;
data_ina = 16'hff26;
data_inb = 16'hffcb;
#10;
address_ina = 78;
address_inb = 79;
data_ina = 16'hf9f0;
data_inb = 16'h3dd;
#10;
address_ina = 80;
address_inb = 81;
data_ina = 16'hff50;
data_inb = 16'hfdaf;
#10;
address_ina = 82;
address_inb = 83;
data_ina = 16'h13f;
data_inb = 16'h570;
#10;
address_ina = 84;
address_inb = 85;
data_ina = 16'h3b6;
data_inb = 16'hff94;
#10;
address_ina = 86;
address_inb = 87;
data_ina = 16'h555;
data_inb = 16'hfdc4;
#10;
address_ina = 88;
address_inb = 89;
data_ina = 16'h1ea;
data_inb = 16'h628;
#10;
address_ina = 90;
address_inb = 91;
data_ina = 16'h596;
data_inb = 16'h38a;
#10;
address_ina = 92;
address_inb = 93;
data_ina = 16'hfbeb;
data_inb = 16'h221;
#10;
address_ina = 94;
address_inb = 95;
data_ina = 16'h36f;
data_inb = 16'hfc2d;
#10;
address_ina = 96;
address_inb = 97;
data_ina = 16'hfdc2;
data_inb = 16'h0;
#10;
address_ina = 98;
address_inb = 99;
data_ina = 16'hfb97;
data_inb = 16'hfe15;
#10;
address_ina = 100;
address_inb = 101;
data_ina = 16'hfed5;
data_inb = 16'hfec3;
#10;
address_ina = 102;
address_inb = 103;
data_ina = 16'h161;
data_inb = 16'hf9f7;
#10;
address_ina = 104;
address_inb = 105;
data_ina = 16'h428;
data_inb = 16'h244;
#10;
address_ina = 106;
address_inb = 107;
data_ina = 16'hf9e4;
data_inb = 16'hff36;
#10;
address_ina = 108;
address_inb = 109;
data_ina = 16'h2dd;
data_inb = 16'hffa0;
#10;
address_ina = 110;
address_inb = 111;
data_ina = 16'h166;
data_inb = 16'hfdd4;
#10;
address_ina = 112;
address_inb = 113;
data_ina = 16'hfe77;
data_inb = 16'h277;
#10;
address_ina = 114;
address_inb = 115;
data_ina = 16'h449;
data_inb = 16'hfdc1;
#10;
address_ina = 116;
address_inb = 117;
data_ina = 16'h4b1;
data_inb = 16'hfcf7;
#10;
address_ina = 118;
address_inb = 119;
data_ina = 16'hfc2d;
data_inb = 16'hd4;
#10;
address_ina = 120;
address_inb = 121;
data_ina = 16'hfc92;
data_inb = 16'hff88;
#10;
address_ina = 122;
address_inb = 123;
data_ina = 16'hfc76;
data_inb = 16'h512;
#10;
address_ina = 124;
address_inb = 125;
data_ina = 16'h62e;
data_inb = 16'hffa2;
#10;
address_ina = 126;
address_inb = 127;
data_ina = 16'h78;
data_inb = 16'hfc58;
#10;
address_ina = 128;
address_inb = 129;
data_ina = 16'hfc65;
data_inb = 16'h63;
#10;
address_ina = 130;
address_inb = 131;
data_ina = 16'h8b;
data_inb = 16'h29;
#10;
address_ina = 132;
address_inb = 133;
data_ina = 16'h33b;
data_inb = 16'h48b;
#10;
address_ina = 134;
address_inb = 135;
data_ina = 16'h518;
data_inb = 16'h5eb;
#10;
address_ina = 136;
address_inb = 137;
data_ina = 16'hfe46;
data_inb = 16'hfa10;
#10;
address_ina = 138;
address_inb = 139;
data_ina = 16'h18a;
data_inb = 16'hfdf9;
#10;
address_ina = 140;
address_inb = 141;
data_ina = 16'hab;
data_inb = 16'hffde;
#10;
address_ina = 142;
address_inb = 143;
data_ina = 16'h5d0;
data_inb = 16'h321;
#10;
address_ina = 144;
address_inb = 145;
data_ina = 16'hfd0b;
data_inb = 16'h29;
#10;
address_ina = 146;
address_inb = 147;
data_ina = 16'h2a6;
data_inb = 16'h3ca;
#10;
address_ina = 148;
address_inb = 149;
data_ina = 16'h5;
data_inb = 16'h397;
#10;
address_ina = 150;
address_inb = 151;
data_ina = 16'hfcfa;
data_inb = 16'h1ee;
#10;
address_ina = 152;
address_inb = 153;
data_ina = 16'hff90;
data_inb = 16'hfc5e;
#10;
address_ina = 154;
address_inb = 155;
data_ina = 16'h2d8;
data_inb = 16'h18e;
#10;
address_ina = 156;
address_inb = 157;
data_ina = 16'h3d0;
data_inb = 16'hfd90;
#10;
address_ina = 158;
address_inb = 159;
data_ina = 16'hfb93;
data_inb = 16'hffe3;
#10;
address_ina = 160;
address_inb = 161;
data_ina = 16'h664;
data_inb = 16'h654;
#10;
address_ina = 162;
address_inb = 163;
data_ina = 16'hfd4d;
data_inb = 16'h2a5;
#10;
address_ina = 164;
address_inb = 165;
data_ina = 16'h3c;
data_inb = 16'hfd76;
#10;
address_ina = 166;
address_inb = 167;
data_ina = 16'hfad4;
data_inb = 16'h108;
#10;
address_ina = 168;
address_inb = 169;
data_ina = 16'h423;
data_inb = 16'h50d;
#10;
address_ina = 170;
address_inb = 171;
data_ina = 16'hfce2;
data_inb = 16'h4c4;
#10;
address_ina = 172;
address_inb = 173;
data_ina = 16'hfa75;
data_inb = 16'h2b5;
#10;
address_ina = 174;
address_inb = 175;
data_ina = 16'h59d;
data_inb = 16'h406;
#10;
address_ina = 176;
address_inb = 177;
data_ina = 16'h529;
data_inb = 16'h5de;
#10;
address_ina = 178;
address_inb = 179;
data_ina = 16'h28a;
data_inb = 16'h25b;
#10;
address_ina = 180;
address_inb = 181;
data_ina = 16'hfd80;
data_inb = 16'h614;
#10;
address_ina = 182;
address_inb = 183;
data_ina = 16'h229;
data_inb = 16'h637;
#10;
address_ina = 184;
address_inb = 185;
data_ina = 16'hf9ad;
data_inb = 16'hfc55;
#10;
address_ina = 186;
address_inb = 187;
data_ina = 16'hfabc;
data_inb = 16'hffe9;
#10;
address_ina = 188;
address_inb = 189;
data_ina = 16'hfb69;
data_inb = 16'h3f2;
#10;
address_ina = 190;
address_inb = 191;
data_ina = 16'h1b2;
data_inb = 16'h508;
#10;
address_ina = 192;
address_inb = 193;
data_ina = 16'hff0f;
data_inb = 16'hfc9f;
#10;
address_ina = 194;
address_inb = 195;
data_ina = 16'h232;
data_inb = 16'h225;
#10;
address_ina = 196;
address_inb = 197;
data_ina = 16'hfe6b;
data_inb = 16'h111;
#10;
address_ina = 198;
address_inb = 199;
data_ina = 16'h3e7;
data_inb = 16'h627;
#10;
address_ina = 200;
address_inb = 201;
data_ina = 16'h15;
data_inb = 16'h167;
#10;
address_ina = 202;
address_inb = 203;
data_ina = 16'h486;
data_inb = 16'hfbeb;
#10;
address_ina = 204;
address_inb = 205;
data_ina = 16'hfeda;
data_inb = 16'h3c6;
#10;
address_ina = 206;
address_inb = 207;
data_ina = 16'hfe10;
data_inb = 16'h1e4;
#10;
address_ina = 208;
address_inb = 209;
data_ina = 16'hff30;
data_inb = 16'h128;
#10;
address_ina = 210;
address_inb = 211;
data_ina = 16'hfdf9;
data_inb = 16'h3b0;
#10;
address_ina = 212;
address_inb = 213;
data_ina = 16'hfbc4;
data_inb = 16'h3c3;
#10;
address_ina = 214;
address_inb = 215;
data_ina = 16'hfed7;
data_inb = 16'h11f;
#10;
address_ina = 216;
address_inb = 217;
data_ina = 16'hb2;
data_inb = 16'h25a;
#10;
address_ina = 218;
address_inb = 219;
data_ina = 16'h3f1;
data_inb = 16'h28c;
#10;
address_ina = 220;
address_inb = 221;
data_ina = 16'hfcea;
data_inb = 16'hfaeb;
#10;
address_ina = 222;
address_inb = 223;
data_ina = 16'h210;
data_inb = 16'hffe0;
#10;
address_ina = 224;
address_inb = 225;
data_ina = 16'hfbd9;
data_inb = 16'hfc1e;
#10;
address_ina = 226;
address_inb = 227;
data_ina = 16'h55d;
data_inb = 16'h3fb;
#10;
address_ina = 228;
address_inb = 229;
data_ina = 16'hfeb6;
data_inb = 16'hff49;
#10;
address_ina = 230;
address_inb = 231;
data_ina = 16'h84;
data_inb = 16'h468;
#10;
address_ina = 232;
address_inb = 233;
data_ina = 16'h310;
data_inb = 16'hfe56;
#10;
address_ina = 234;
address_inb = 235;
data_ina = 16'hffd2;
data_inb = 16'h47e;
#10;
address_ina = 236;
address_inb = 237;
data_ina = 16'h36b;
data_inb = 16'h30c;
#10;
address_ina = 238;
address_inb = 239;
data_ina = 16'h1d9;
data_inb = 16'h1bb;
#10;
address_ina = 240;
address_inb = 241;
data_ina = 16'hfea0;
data_inb = 16'h23e;
#10;
address_ina = 242;
address_inb = 243;
data_ina = 16'hfb20;
data_inb = 16'hfd2a;
#10;
address_ina = 244;
address_inb = 245;
data_ina = 16'hfd81;
data_inb = 16'h142;
#10;
address_ina = 246;
address_inb = 247;
data_ina = 16'h263;
data_inb = 16'hff16;
#10;
address_ina = 248;
address_inb = 249;
data_ina = 16'hfc54;
data_inb = 16'h188;
#10;
address_ina = 250;
address_inb = 251;
data_ina = 16'hfa71;
data_inb = 16'hfd96;
#10;
address_ina = 252;
address_inb = 253;
data_ina = 16'h48a;
data_inb = 16'hfe00;
#10;
address_ina = 254;
address_inb = 255;
data_ina = 16'h5cc;
data_inb = 16'h7a;
#10;
        wait(init_done);
        #30
        we = 0;
        // Start processing
         
		  #38000

        start = 0;



//        wait (wr_req);
//		  wait (!wr_req);
//		   rd_req = 1;
		  wait(done);
		  #20000
rd_req = 1;
        #70 
		  start = 1;
		 #80 
wait(rd_empty)
rd_req = 0;

$display("Finished the NTT test Number %d",test_num);
////Begin test number #100//////////////
rst = 1;

//#1000
start = 1;
mode = 1; //NTT 0 // INTT 1

// Reset for a few clock cycles

#1000

rst = 0;
test_num = test_num + 1;
#1000
we = 1;
address_ina = 0;
address_inb = 1;
data_ina = 16'hfc85;
data_inb = 16'h664;
#10;
address_ina = 2;
address_inb = 3;
data_ina = 16'hfa0d;
data_inb = 16'h60f;
#10;
address_ina = 4;
address_inb = 5;
data_ina = 16'hff0c;
data_inb = 16'hfa28;
#10;
address_ina = 6;
address_inb = 7;
data_ina = 16'h90;
data_inb = 16'h18e;
#10;
address_ina = 8;
address_inb = 9;
data_ina = 16'h4fc;
data_inb = 16'hfaee;
#10;
address_ina = 10;
address_inb = 11;
data_ina = 16'h677;
data_inb = 16'h463;
#10;
address_ina = 12;
address_inb = 13;
data_ina = 16'h433;
data_inb = 16'hfc0d;
#10;
address_ina = 14;
address_inb = 15;
data_ina = 16'hd5;
data_inb = 16'hfec0;
#10;
address_ina = 16;
address_inb = 17;
data_ina = 16'hfe23;
data_inb = 16'h53c;
#10;
address_ina = 18;
address_inb = 19;
data_ina = 16'h149;
data_inb = 16'h4ed;
#10;
address_ina = 20;
address_inb = 21;
data_ina = 16'h67a;
data_inb = 16'hff0a;
#10;
address_ina = 22;
address_inb = 23;
data_ina = 16'h3f6;
data_inb = 16'hff52;
#10;
address_ina = 24;
address_inb = 25;
data_ina = 16'hfce3;
data_inb = 16'hfc70;
#10;
address_ina = 26;
address_inb = 27;
data_ina = 16'h82;
data_inb = 16'hfc47;
#10;
address_ina = 28;
address_inb = 29;
data_ina = 16'hfa6d;
data_inb = 16'h29e;
#10;
address_ina = 30;
address_inb = 31;
data_ina = 16'hfc76;
data_inb = 16'h59b;
#10;
address_ina = 32;
address_inb = 33;
data_ina = 16'hffff;
data_inb = 16'hfdce;
#10;
address_ina = 34;
address_inb = 35;
data_ina = 16'h1d4;
data_inb = 16'hfbbe;
#10;
address_ina = 36;
address_inb = 37;
data_ina = 16'h5b6;
data_inb = 16'hfe64;
#10;
address_ina = 38;
address_inb = 39;
data_ina = 16'h629;
data_inb = 16'h28a;
#10;
address_ina = 40;
address_inb = 41;
data_ina = 16'hfe0d;
data_inb = 16'hfe64;
#10;
address_ina = 42;
address_inb = 43;
data_ina = 16'h31c;
data_inb = 16'hfd41;
#10;
address_ina = 44;
address_inb = 45;
data_ina = 16'hffd0;
data_inb = 16'h48a;
#10;
address_ina = 46;
address_inb = 47;
data_ina = 16'hfba2;
data_inb = 16'hb6;
#10;
address_ina = 48;
address_inb = 49;
data_ina = 16'h332;
data_inb = 16'h0;
#10;
address_ina = 50;
address_inb = 51;
data_ina = 16'h572;
data_inb = 16'h4ed;
#10;
address_ina = 52;
address_inb = 53;
data_ina = 16'h3d;
data_inb = 16'hfe90;
#10;
address_ina = 54;
address_inb = 55;
data_ina = 16'hf989;
data_inb = 16'hfe03;
#10;
address_ina = 56;
address_inb = 57;
data_ina = 16'h1c0;
data_inb = 16'h382;
#10;
address_ina = 58;
address_inb = 59;
data_ina = 16'hfec2;
data_inb = 16'h5b1;
#10;
address_ina = 60;
address_inb = 61;
data_ina = 16'hfd7d;
data_inb = 16'h3ec;
#10;
address_ina = 62;
address_inb = 63;
data_ina = 16'hfb20;
data_inb = 16'hfc92;
#10;
address_ina = 64;
address_inb = 65;
data_ina = 16'hfc06;
data_inb = 16'h4dd;
#10;
address_ina = 66;
address_inb = 67;
data_ina = 16'h315;
data_inb = 16'h1cf;
#10;
address_ina = 68;
address_inb = 69;
data_ina = 16'h192;
data_inb = 16'h2c0;
#10;
address_ina = 70;
address_inb = 71;
data_ina = 16'hfffe;
data_inb = 16'hff34;
#10;
address_ina = 72;
address_inb = 73;
data_ina = 16'hff00;
data_inb = 16'hfcb5;
#10;
address_ina = 74;
address_inb = 75;
data_ina = 16'hfa0c;
data_inb = 16'h5ec;
#10;
address_ina = 76;
address_inb = 77;
data_ina = 16'hfc19;
data_inb = 16'h5f3;
#10;
address_ina = 78;
address_inb = 79;
data_ina = 16'h4fe;
data_inb = 16'h19b;
#10;
address_ina = 80;
address_inb = 81;
data_ina = 16'hfad4;
data_inb = 16'h1f3;
#10;
address_ina = 82;
address_inb = 83;
data_ina = 16'h482;
data_inb = 16'hfc27;
#10;
address_ina = 84;
address_inb = 85;
data_ina = 16'hfa8d;
data_inb = 16'hfb4e;
#10;
address_ina = 86;
address_inb = 87;
data_ina = 16'h31e;
data_inb = 16'hfb23;
#10;
address_ina = 88;
address_inb = 89;
data_ina = 16'h2f4;
data_inb = 16'h11e;
#10;
address_ina = 90;
address_inb = 91;
data_ina = 16'hfde6;
data_inb = 16'h5d4;
#10;
address_ina = 92;
address_inb = 93;
data_ina = 16'hfc14;
data_inb = 16'hfdbd;
#10;
address_ina = 94;
address_inb = 95;
data_ina = 16'h294;
data_inb = 16'h2b4;
#10;
address_ina = 96;
address_inb = 97;
data_ina = 16'h138;
data_inb = 16'h42d;
#10;
address_ina = 98;
address_inb = 99;
data_ina = 16'hfd5f;
data_inb = 16'hffa8;
#10;
address_ina = 100;
address_inb = 101;
data_ina = 16'h113;
data_inb = 16'h28d;
#10;
address_ina = 102;
address_inb = 103;
data_ina = 16'h320;
data_inb = 16'h52f;
#10;
address_ina = 104;
address_inb = 105;
data_ina = 16'h645;
data_inb = 16'hfeb4;
#10;
address_ina = 106;
address_inb = 107;
data_ina = 16'h118;
data_inb = 16'hfb69;
#10;
address_ina = 108;
address_inb = 109;
data_ina = 16'hfe59;
data_inb = 16'hfd33;
#10;
address_ina = 110;
address_inb = 111;
data_ina = 16'hc;
data_inb = 16'hfbcf;
#10;
address_ina = 112;
address_inb = 113;
data_ina = 16'h46;
data_inb = 16'hff10;
#10;
address_ina = 114;
address_inb = 115;
data_ina = 16'hfdc8;
data_inb = 16'hfbdf;
#10;
address_ina = 116;
address_inb = 117;
data_ina = 16'h49e;
data_inb = 16'hfec2;
#10;
address_ina = 118;
address_inb = 119;
data_ina = 16'hfba8;
data_inb = 16'hfff3;
#10;
address_ina = 120;
address_inb = 121;
data_ina = 16'h35f;
data_inb = 16'hfebb;
#10;
address_ina = 122;
address_inb = 123;
data_ina = 16'hff25;
data_inb = 16'h503;
#10;
address_ina = 124;
address_inb = 125;
data_ina = 16'hfb07;
data_inb = 16'hfbab;
#10;
address_ina = 126;
address_inb = 127;
data_ina = 16'h1fe;
data_inb = 16'h7d;
#10;
address_ina = 128;
address_inb = 129;
data_ina = 16'hfa74;
data_inb = 16'h5eb;
#10;
address_ina = 130;
address_inb = 131;
data_ina = 16'hff6d;
data_inb = 16'h312;
#10;
address_ina = 132;
address_inb = 133;
data_ina = 16'h3ea;
data_inb = 16'hfcb9;
#10;
address_ina = 134;
address_inb = 135;
data_ina = 16'hfb91;
data_inb = 16'hfb43;
#10;
address_ina = 136;
address_inb = 137;
data_ina = 16'hf9ab;
data_inb = 16'hfba9;
#10;
address_ina = 138;
address_inb = 139;
data_ina = 16'hfc92;
data_inb = 16'h222;
#10;
address_ina = 140;
address_inb = 141;
data_ina = 16'hec;
data_inb = 16'hff14;
#10;
address_ina = 142;
address_inb = 143;
data_ina = 16'h2c1;
data_inb = 16'hfa5e;
#10;
address_ina = 144;
address_inb = 145;
data_ina = 16'h177;
data_inb = 16'hfbfc;
#10;
address_ina = 146;
address_inb = 147;
data_ina = 16'h3a;
data_inb = 16'hfbc8;
#10;
address_ina = 148;
address_inb = 149;
data_ina = 16'h102;
data_inb = 16'hfb7f;
#10;
address_ina = 150;
address_inb = 151;
data_ina = 16'h2a8;
data_inb = 16'hfc32;
#10;
address_ina = 152;
address_inb = 153;
data_ina = 16'hfda2;
data_inb = 16'hfdee;
#10;
address_ina = 154;
address_inb = 155;
data_ina = 16'hfbb4;
data_inb = 16'h385;
#10;
address_ina = 156;
address_inb = 157;
data_ina = 16'h561;
data_inb = 16'hfeab;
#10;
address_ina = 158;
address_inb = 159;
data_ina = 16'hfeef;
data_inb = 16'hfcf0;
#10;
address_ina = 160;
address_inb = 161;
data_ina = 16'h57f;
data_inb = 16'h66;
#10;
address_ina = 162;
address_inb = 163;
data_ina = 16'hfd0b;
data_inb = 16'h1af;
#10;
address_ina = 164;
address_inb = 165;
data_ina = 16'hfec0;
data_inb = 16'hfec5;
#10;
address_ina = 166;
address_inb = 167;
data_ina = 16'h2ed;
data_inb = 16'hf9f1;
#10;
address_ina = 168;
address_inb = 169;
data_ina = 16'h119;
data_inb = 16'h21;
#10;
address_ina = 170;
address_inb = 171;
data_ina = 16'h21b;
data_inb = 16'h411;
#10;
address_ina = 172;
address_inb = 173;
data_ina = 16'h3a9;
data_inb = 16'hfe4f;
#10;
address_ina = 174;
address_inb = 175;
data_ina = 16'hffeb;
data_inb = 16'hfe4f;
#10;
address_ina = 176;
address_inb = 177;
data_ina = 16'h2fd;
data_inb = 16'hf9a6;
#10;
address_ina = 178;
address_inb = 179;
data_ina = 16'hff9d;
data_inb = 16'hfc82;
#10;
address_ina = 180;
address_inb = 181;
data_ina = 16'h2a;
data_inb = 16'hfc5d;
#10;
address_ina = 182;
address_inb = 183;
data_ina = 16'hfb94;
data_inb = 16'h4a0;
#10;
address_ina = 184;
address_inb = 185;
data_ina = 16'hfc9e;
data_inb = 16'hfe00;
#10;
address_ina = 186;
address_inb = 187;
data_ina = 16'hfa70;
data_inb = 16'hfc7b;
#10;
address_ina = 188;
address_inb = 189;
data_ina = 16'hfd41;
data_inb = 16'h452;
#10;
address_ina = 190;
address_inb = 191;
data_ina = 16'h537;
data_inb = 16'h3c6;
#10;
address_ina = 192;
address_inb = 193;
data_ina = 16'hfa45;
data_inb = 16'hff18;
#10;
address_ina = 194;
address_inb = 195;
data_ina = 16'hfde1;
data_inb = 16'hffa2;
#10;
address_ina = 196;
address_inb = 197;
data_ina = 16'h31f;
data_inb = 16'hfdf8;
#10;
address_ina = 198;
address_inb = 199;
data_ina = 16'h678;
data_inb = 16'h636;
#10;
address_ina = 200;
address_inb = 201;
data_ina = 16'h344;
data_inb = 16'hffa8;
#10;
address_ina = 202;
address_inb = 203;
data_ina = 16'hfde1;
data_inb = 16'hfa4e;
#10;
address_ina = 204;
address_inb = 205;
data_ina = 16'h5ab;
data_inb = 16'h40c;
#10;
address_ina = 206;
address_inb = 207;
data_ina = 16'hf9a5;
data_inb = 16'h1e1;
#10;
address_ina = 208;
address_inb = 209;
data_ina = 16'hf9f0;
data_inb = 16'h1cc;
#10;
address_ina = 210;
address_inb = 211;
data_ina = 16'hfe10;
data_inb = 16'h315;
#10;
address_ina = 212;
address_inb = 213;
data_ina = 16'h1e7;
data_inb = 16'h20e;
#10;
address_ina = 214;
address_inb = 215;
data_ina = 16'h648;
data_inb = 16'hfc69;
#10;
address_ina = 216;
address_inb = 217;
data_ina = 16'hff5a;
data_inb = 16'he7;
#10;
address_ina = 218;
address_inb = 219;
data_ina = 16'hfa43;
data_inb = 16'h4d2;
#10;
address_ina = 220;
address_inb = 221;
data_ina = 16'hfd43;
data_inb = 16'h352;
#10;
address_ina = 222;
address_inb = 223;
data_ina = 16'h15e;
data_inb = 16'hf9bf;
#10;
address_ina = 224;
address_inb = 225;
data_ina = 16'hff96;
data_inb = 16'hfc64;
#10;
address_ina = 226;
address_inb = 227;
data_ina = 16'hfbfa;
data_inb = 16'h6f;
#10;
address_ina = 228;
address_inb = 229;
data_ina = 16'h1e0;
data_inb = 16'hf98d;
#10;
address_ina = 230;
address_inb = 231;
data_ina = 16'h580;
data_inb = 16'hfb49;
#10;
address_ina = 232;
address_inb = 233;
data_ina = 16'h669;
data_inb = 16'hfd8c;
#10;
address_ina = 234;
address_inb = 235;
data_ina = 16'hfb29;
data_inb = 16'hff9f;
#10;
address_ina = 236;
address_inb = 237;
data_ina = 16'h46b;
data_inb = 16'hff9f;
#10;
address_ina = 238;
address_inb = 239;
data_ina = 16'h5a1;
data_inb = 16'hff37;
#10;
address_ina = 240;
address_inb = 241;
data_ina = 16'h120;
data_inb = 16'h28a;
#10;
address_ina = 242;
address_inb = 243;
data_ina = 16'h74;
data_inb = 16'h3a9;
#10;
address_ina = 244;
address_inb = 245;
data_ina = 16'h64;
data_inb = 16'h370;
#10;
address_ina = 246;
address_inb = 247;
data_ina = 16'h5f;
data_inb = 16'hf985;
#10;
address_ina = 248;
address_inb = 249;
data_ina = 16'h434;
data_inb = 16'h3ed;
#10;
address_ina = 250;
address_inb = 251;
data_ina = 16'h5e6;
data_inb = 16'h2dc;
#10;
address_ina = 252;
address_inb = 253;
data_ina = 16'hfe60;
data_inb = 16'h56a;
#10;
address_ina = 254;
address_inb = 255;
data_ina = 16'h402;
data_inb = 16'h20f;
#10;
        wait(init_done);
        #30
        we = 0;
        // Start processing
         
		  #38000

        start = 0;



//        wait (wr_req);
//		  wait (!wr_req);
//		   rd_req = 1;
		  wait(done);
		  #20000
rd_req = 1;
        #70 
		  start = 1;
		 #80 
wait(rd_empty)
rd_req = 0;

$display("Finished the NTT test Number %d",test_num);
////Begin test number #101//////////////
rst = 1;

//#1000
start = 1;
mode = 1; //NTT 0 // INTT 1

// Reset for a few clock cycles

#1000

rst = 0;
test_num = test_num + 1;
#1000
we = 1;
address_ina = 0;
address_inb = 1;
data_ina = 16'hfd10;
data_inb = 16'hfd43;
#10;
address_ina = 2;
address_inb = 3;
data_ina = 16'h6a;
data_inb = 16'hf9fa;
#10;
address_ina = 4;
address_inb = 5;
data_ina = 16'hfba4;
data_inb = 16'hfb53;
#10;
address_ina = 6;
address_inb = 7;
data_ina = 16'h394;
data_inb = 16'hfa0b;
#10;
address_ina = 8;
address_inb = 9;
data_ina = 16'h30;
data_inb = 16'h667;
#10;
address_ina = 10;
address_inb = 11;
data_ina = 16'hfd36;
data_inb = 16'hfaa4;
#10;
address_ina = 12;
address_inb = 13;
data_ina = 16'hf9ce;
data_inb = 16'h32e;
#10;
address_ina = 14;
address_inb = 15;
data_ina = 16'h3c5;
data_inb = 16'hfe61;
#10;
address_ina = 16;
address_inb = 17;
data_ina = 16'hfe99;
data_inb = 16'h345;
#10;
address_ina = 18;
address_inb = 19;
data_ina = 16'h26e;
data_inb = 16'hfd70;
#10;
address_ina = 20;
address_inb = 21;
data_ina = 16'h180;
data_inb = 16'hfa75;
#10;
address_ina = 22;
address_inb = 23;
data_ina = 16'h1ec;
data_inb = 16'h199;
#10;
address_ina = 24;
address_inb = 25;
data_ina = 16'h3df;
data_inb = 16'h3f3;
#10;
address_ina = 26;
address_inb = 27;
data_ina = 16'hfbc4;
data_inb = 16'h46a;
#10;
address_ina = 28;
address_inb = 29;
data_ina = 16'h59d;
data_inb = 16'hff00;
#10;
address_ina = 30;
address_inb = 31;
data_ina = 16'hf9b5;
data_inb = 16'hfabc;
#10;
address_ina = 32;
address_inb = 33;
data_ina = 16'h40d;
data_inb = 16'h566;
#10;
address_ina = 34;
address_inb = 35;
data_ina = 16'hfdd9;
data_inb = 16'h4;
#10;
address_ina = 36;
address_inb = 37;
data_ina = 16'hffad;
data_inb = 16'hbd;
#10;
address_ina = 38;
address_inb = 39;
data_ina = 16'hfe0d;
data_inb = 16'h1ca;
#10;
address_ina = 40;
address_inb = 41;
data_ina = 16'hfc13;
data_inb = 16'h62b;
#10;
address_ina = 42;
address_inb = 43;
data_ina = 16'h5b2;
data_inb = 16'h275;
#10;
address_ina = 44;
address_inb = 45;
data_ina = 16'hf9b3;
data_inb = 16'hff0e;
#10;
address_ina = 46;
address_inb = 47;
data_ina = 16'hff75;
data_inb = 16'h91;
#10;
address_ina = 48;
address_inb = 49;
data_ina = 16'hfb33;
data_inb = 16'h18c;
#10;
address_ina = 50;
address_inb = 51;
data_ina = 16'h35;
data_inb = 16'h11c;
#10;
address_ina = 52;
address_inb = 53;
data_ina = 16'hfe8d;
data_inb = 16'hfade;
#10;
address_ina = 54;
address_inb = 55;
data_ina = 16'hf99e;
data_inb = 16'h603;
#10;
address_ina = 56;
address_inb = 57;
data_ina = 16'h82;
data_inb = 16'h18e;
#10;
address_ina = 58;
address_inb = 59;
data_ina = 16'h454;
data_inb = 16'hfe72;
#10;
address_ina = 60;
address_inb = 61;
data_ina = 16'h5b2;
data_inb = 16'h407;
#10;
address_ina = 62;
address_inb = 63;
data_ina = 16'h647;
data_inb = 16'hfd54;
#10;
address_ina = 64;
address_inb = 65;
data_ina = 16'h1a6;
data_inb = 16'hfe1e;
#10;
address_ina = 66;
address_inb = 67;
data_ina = 16'h439;
data_inb = 16'h45f;
#10;
address_ina = 68;
address_inb = 69;
data_ina = 16'h353;
data_inb = 16'h4c0;
#10;
address_ina = 70;
address_inb = 71;
data_ina = 16'hf9d5;
data_inb = 16'h424;
#10;
address_ina = 72;
address_inb = 73;
data_ina = 16'hfc8d;
data_inb = 16'hff7c;
#10;
address_ina = 74;
address_inb = 75;
data_ina = 16'h194;
data_inb = 16'h10f;
#10;
address_ina = 76;
address_inb = 77;
data_ina = 16'hd7;
data_inb = 16'h10b;
#10;
address_ina = 78;
address_inb = 79;
data_ina = 16'hfb0b;
data_inb = 16'hfd13;
#10;
address_ina = 80;
address_inb = 81;
data_ina = 16'hec;
data_inb = 16'hfc09;
#10;
address_ina = 82;
address_inb = 83;
data_ina = 16'hfd6a;
data_inb = 16'h5c3;
#10;
address_ina = 84;
address_inb = 85;
data_ina = 16'hfaa2;
data_inb = 16'h384;
#10;
address_ina = 86;
address_inb = 87;
data_ina = 16'h36d;
data_inb = 16'h5a9;
#10;
address_ina = 88;
address_inb = 89;
data_ina = 16'hfb56;
data_inb = 16'hfcce;
#10;
address_ina = 90;
address_inb = 91;
data_ina = 16'h74;
data_inb = 16'hfb17;
#10;
address_ina = 92;
address_inb = 93;
data_ina = 16'h5da;
data_inb = 16'hfdbc;
#10;
address_ina = 94;
address_inb = 95;
data_ina = 16'h459;
data_inb = 16'he0;
#10;
address_ina = 96;
address_inb = 97;
data_ina = 16'h5b4;
data_inb = 16'hfef4;
#10;
address_ina = 98;
address_inb = 99;
data_ina = 16'h54d;
data_inb = 16'h5d7;
#10;
address_ina = 100;
address_inb = 101;
data_ina = 16'h188;
data_inb = 16'h35c;
#10;
address_ina = 102;
address_inb = 103;
data_ina = 16'hfa7f;
data_inb = 16'hfd56;
#10;
address_ina = 104;
address_inb = 105;
data_ina = 16'hfed2;
data_inb = 16'h4;
#10;
address_ina = 106;
address_inb = 107;
data_ina = 16'hfe52;
data_inb = 16'h2ff;
#10;
address_ina = 108;
address_inb = 109;
data_ina = 16'h268;
data_inb = 16'h23b;
#10;
address_ina = 110;
address_inb = 111;
data_ina = 16'h407;
data_inb = 16'hfae9;
#10;
address_ina = 112;
address_inb = 113;
data_ina = 16'h9e;
data_inb = 16'h3b7;
#10;
address_ina = 114;
address_inb = 115;
data_ina = 16'hfd1c;
data_inb = 16'hfc09;
#10;
address_ina = 116;
address_inb = 117;
data_ina = 16'h234;
data_inb = 16'h62e;
#10;
address_ina = 118;
address_inb = 119;
data_ina = 16'hfb3b;
data_inb = 16'hfd4a;
#10;
address_ina = 120;
address_inb = 121;
data_ina = 16'hfae6;
data_inb = 16'h4fe;
#10;
address_ina = 122;
address_inb = 123;
data_ina = 16'h261;
data_inb = 16'h528;
#10;
address_ina = 124;
address_inb = 125;
data_ina = 16'h19e;
data_inb = 16'h2f9;
#10;
address_ina = 126;
address_inb = 127;
data_ina = 16'hfbf8;
data_inb = 16'hfe98;
#10;
address_ina = 128;
address_inb = 129;
data_ina = 16'h19e;
data_inb = 16'h230;
#10;
address_ina = 130;
address_inb = 131;
data_ina = 16'hcb;
data_inb = 16'h3d2;
#10;
address_ina = 132;
address_inb = 133;
data_ina = 16'hfa46;
data_inb = 16'h135;
#10;
address_ina = 134;
address_inb = 135;
data_ina = 16'h1b5;
data_inb = 16'hd;
#10;
address_ina = 136;
address_inb = 137;
data_ina = 16'h60b;
data_inb = 16'hfec9;
#10;
address_ina = 138;
address_inb = 139;
data_ina = 16'h3;
data_inb = 16'h2bd;
#10;
address_ina = 140;
address_inb = 141;
data_ina = 16'hfe4c;
data_inb = 16'hfca2;
#10;
address_ina = 142;
address_inb = 143;
data_ina = 16'h2a;
data_inb = 16'h248;
#10;
address_ina = 144;
address_inb = 145;
data_ina = 16'hfb88;
data_inb = 16'hfae5;
#10;
address_ina = 146;
address_inb = 147;
data_ina = 16'hfece;
data_inb = 16'hfea1;
#10;
address_ina = 148;
address_inb = 149;
data_ina = 16'hfda8;
data_inb = 16'hf999;
#10;
address_ina = 150;
address_inb = 151;
data_ina = 16'hf994;
data_inb = 16'h3ff;
#10;
address_ina = 152;
address_inb = 153;
data_ina = 16'h8b;
data_inb = 16'h21b;
#10;
address_ina = 154;
address_inb = 155;
data_ina = 16'hfa56;
data_inb = 16'h3af;
#10;
address_ina = 156;
address_inb = 157;
data_ina = 16'h442;
data_inb = 16'hfe28;
#10;
address_ina = 158;
address_inb = 159;
data_ina = 16'hff9c;
data_inb = 16'h666;
#10;
address_ina = 160;
address_inb = 161;
data_ina = 16'h1ec;
data_inb = 16'h292;
#10;
address_ina = 162;
address_inb = 163;
data_ina = 16'h2cb;
data_inb = 16'hfd3a;
#10;
address_ina = 164;
address_inb = 165;
data_ina = 16'hfa62;
data_inb = 16'hffe3;
#10;
address_ina = 166;
address_inb = 167;
data_ina = 16'h52;
data_inb = 16'h396;
#10;
address_ina = 168;
address_inb = 169;
data_ina = 16'ha2;
data_inb = 16'hfc73;
#10;
address_ina = 170;
address_inb = 171;
data_ina = 16'h3a1;
data_inb = 16'haf;
#10;
address_ina = 172;
address_inb = 173;
data_ina = 16'hfff5;
data_inb = 16'hfa8e;
#10;
address_ina = 174;
address_inb = 175;
data_ina = 16'hf3;
data_inb = 16'hfbe8;
#10;
address_ina = 176;
address_inb = 177;
data_ina = 16'h1b0;
data_inb = 16'h5b8;
#10;
address_ina = 178;
address_inb = 179;
data_ina = 16'hfe29;
data_inb = 16'h112;
#10;
address_ina = 180;
address_inb = 181;
data_ina = 16'h286;
data_inb = 16'h567;
#10;
address_ina = 182;
address_inb = 183;
data_ina = 16'h3ca;
data_inb = 16'hfecc;
#10;
address_ina = 184;
address_inb = 185;
data_ina = 16'hff28;
data_inb = 16'hfe00;
#10;
address_ina = 186;
address_inb = 187;
data_ina = 16'hfc8e;
data_inb = 16'hfcd7;
#10;
address_ina = 188;
address_inb = 189;
data_ina = 16'h18f;
data_inb = 16'h2b2;
#10;
address_ina = 190;
address_inb = 191;
data_ina = 16'hf9f8;
data_inb = 16'h61;
#10;
address_ina = 192;
address_inb = 193;
data_ina = 16'hfbd9;
data_inb = 16'h24b;
#10;
address_ina = 194;
address_inb = 195;
data_ina = 16'h5a1;
data_inb = 16'h3f8;
#10;
address_ina = 196;
address_inb = 197;
data_ina = 16'hffbb;
data_inb = 16'hfde6;
#10;
address_ina = 198;
address_inb = 199;
data_ina = 16'hfac8;
data_inb = 16'hfde8;
#10;
address_ina = 200;
address_inb = 201;
data_ina = 16'hfbcf;
data_inb = 16'hfede;
#10;
address_ina = 202;
address_inb = 203;
data_ina = 16'h528;
data_inb = 16'hfe79;
#10;
address_ina = 204;
address_inb = 205;
data_ina = 16'h368;
data_inb = 16'hfbd2;
#10;
address_ina = 206;
address_inb = 207;
data_ina = 16'hfd9c;
data_inb = 16'h665;
#10;
address_ina = 208;
address_inb = 209;
data_ina = 16'hf9ca;
data_inb = 16'hf9dc;
#10;
address_ina = 210;
address_inb = 211;
data_ina = 16'h180;
data_inb = 16'hfcfc;
#10;
address_ina = 212;
address_inb = 213;
data_ina = 16'hfa45;
data_inb = 16'h1fe;
#10;
address_ina = 214;
address_inb = 215;
data_ina = 16'hffb8;
data_inb = 16'h223;
#10;
address_ina = 216;
address_inb = 217;
data_ina = 16'hfd1a;
data_inb = 16'hfdf6;
#10;
address_ina = 218;
address_inb = 219;
data_ina = 16'hfd76;
data_inb = 16'h162;
#10;
address_ina = 220;
address_inb = 221;
data_ina = 16'h25d;
data_inb = 16'h4aa;
#10;
address_ina = 222;
address_inb = 223;
data_ina = 16'h83;
data_inb = 16'h67c;
#10;
address_ina = 224;
address_inb = 225;
data_ina = 16'hfdf8;
data_inb = 16'hfe77;
#10;
address_ina = 226;
address_inb = 227;
data_ina = 16'h283;
data_inb = 16'hfb09;
#10;
address_ina = 228;
address_inb = 229;
data_ina = 16'hfcb0;
data_inb = 16'hfafd;
#10;
address_ina = 230;
address_inb = 231;
data_ina = 16'h25e;
data_inb = 16'h36e;
#10;
address_ina = 232;
address_inb = 233;
data_ina = 16'hfe28;
data_inb = 16'h630;
#10;
address_ina = 234;
address_inb = 235;
data_ina = 16'hfeac;
data_inb = 16'hfe56;
#10;
address_ina = 236;
address_inb = 237;
data_ina = 16'hfa6f;
data_inb = 16'ha2;
#10;
address_ina = 238;
address_inb = 239;
data_ina = 16'h11d;
data_inb = 16'hfb5c;
#10;
address_ina = 240;
address_inb = 241;
data_ina = 16'hb2;
data_inb = 16'h313;
#10;
address_ina = 242;
address_inb = 243;
data_ina = 16'hfbb4;
data_inb = 16'hfaad;
#10;
address_ina = 244;
address_inb = 245;
data_ina = 16'h40c;
data_inb = 16'hf9dd;
#10;
address_ina = 246;
address_inb = 247;
data_ina = 16'h168;
data_inb = 16'hb7;
#10;
address_ina = 248;
address_inb = 249;
data_ina = 16'hfe31;
data_inb = 16'hfb50;
#10;
address_ina = 250;
address_inb = 251;
data_ina = 16'h368;
data_inb = 16'hff80;
#10;
address_ina = 252;
address_inb = 253;
data_ina = 16'h4b6;
data_inb = 16'h117;
#10;
address_ina = 254;
address_inb = 255;
data_ina = 16'h3e;
data_inb = 16'h3fc;
#10;
        wait(init_done);
        #30
        we = 0;
        // Start processing
         
		  #38000

        start = 0;



//        wait (wr_req);
//		  wait (!wr_req);
//		   rd_req = 1;
		  wait(done);
		  #20000
rd_req = 1;
        #70 
		  start = 1;
		 #80 
wait(rd_empty)
rd_req = 0;

$display("Finished the NTT test Number %d",test_num);


$display("Finished all tests");
        $finish; 
    end 

integer filelog;
 
always@(posedge clk)
begin
if(wr_req)
begin
	filelog=$fopen("./log.txt2","a");
    $display("data out 1 = %h ; data out 2 = %h",data_out1,data_out2);
	//$display("data out 2 = %h",data_out2);
	$fwrite(filelog,"current test num = %d, data out 1 = %h ; data out 2 = %h\n",test_num, data_out1, data_out2);
	$fclose(filelog);
end
end

endmodule 

 

 